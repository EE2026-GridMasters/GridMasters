`timescale 1ns / 1ps

module display_mode_select_pvp(
    input [12:0] pixel_index,
    output reg [15:0] oled_data
    );
    
    parameter PINK_HEX = 16'hF899;
    parameter BLUE_HEX = 16'h177F;
    parameter BG_BLUE_HEX = 16'b0000000001000100;
    parameter WHITE_HEX = 16'hFFFF;
    
    always @(*) begin
        if ((pixel_index >= 783 && pixel_index <= 848) || (pixel_index >= 878 && pixel_index <= 945) || (pixel_index >= 973 && pixel_index <= 1042) || (pixel_index >= 1069 && pixel_index <= 1138) || (pixel_index >= 1165 && pixel_index <= 1234) || (pixel_index >= 1261 && pixel_index <= 1276) || (pixel_index >= 1279 && pixel_index <= 1312) || (pixel_index >= 1315 && pixel_index <= 1330) || (pixel_index >= 1357 && pixel_index <= 1372) || (pixel_index >= 1375 && pixel_index <= 1408) || (pixel_index >= 1411 && pixel_index <= 1426) || (pixel_index >= 1453 && pixel_index <= 1464) || (pixel_index >= 1471 && pixel_index <= 1500) || (pixel_index >= 1507 && pixel_index <= 1522) || (pixel_index >= 1549 && pixel_index <= 1560) || (pixel_index >= 1567 && pixel_index <= 1577) || (pixel_index >= 1580 && pixel_index <= 1585) || (pixel_index >= 1588 && pixel_index <= 1596) || (pixel_index >= 1603 && pixel_index <= 1618) || (pixel_index >= 1645 && pixel_index <= 1660) || (pixel_index >= 1663 && pixel_index <= 1673) || (pixel_index >= 1676 && pixel_index <= 1681) || (pixel_index >= 1684 && pixel_index <= 1696) || (pixel_index >= 1699 && pixel_index <= 1714) || (pixel_index >= 1741 && pixel_index <= 1756) || (pixel_index >= 1759 && pixel_index <= 1771) || (pixel_index >= 1774 && pixel_index <= 1775) || (pixel_index >= 1778 && pixel_index <= 1792) || (pixel_index >= 1795 && pixel_index <= 1810) || (pixel_index >= 1837 && pixel_index <= 1852) || (pixel_index >= 1855 && pixel_index <= 1867) || (pixel_index >= 1870 && pixel_index <= 1871) || (pixel_index >= 1874 && pixel_index <= 1888) || (pixel_index >= 1891 && pixel_index <= 1906) || (pixel_index >= 1933 && pixel_index <= 1948) || (pixel_index >= 1951 && pixel_index <= 1963) || (pixel_index >= 1966 && pixel_index <= 1967) || (pixel_index >= 1970 && pixel_index <= 1984) || (pixel_index >= 1987 && pixel_index <= 2002) || (pixel_index >= 2029 && pixel_index <= 2044) || (pixel_index >= 2047 && pixel_index <= 2059) || (pixel_index >= 2062 && pixel_index <= 2063) || (pixel_index >= 2066 && pixel_index <= 2080) || (pixel_index >= 2083 && pixel_index <= 2098) || (pixel_index >= 2125 && pixel_index <= 2140) || (pixel_index >= 2143 && pixel_index <= 2157) || (pixel_index >= 2160 && pixel_index <= 2176) || (pixel_index >= 2179 && pixel_index <= 2194) || (pixel_index >= 2221 && pixel_index <= 2236) || (pixel_index >= 2239 && pixel_index <= 2253) || (pixel_index >= 2256 && pixel_index <= 2272) || (pixel_index >= 2275 && pixel_index <= 2290) || (pixel_index >= 2317 && pixel_index <= 2332) || (pixel_index >= 2335 && pixel_index <= 2349) || (pixel_index >= 2352 && pixel_index <= 2368) || (pixel_index >= 2371 && pixel_index <= 2386) || (pixel_index >= 2413 && pixel_index <= 2428) || (pixel_index >= 2431 && pixel_index <= 2445) || (pixel_index >= 2448 && pixel_index <= 2464) || (pixel_index >= 2467 && pixel_index <= 2482) || (pixel_index >= 2509 && pixel_index <= 2578) || (pixel_index >= 2605 && pixel_index <= 2674) || (pixel_index >= 2701 && pixel_index <= 2770) || (pixel_index >= 2798 && pixel_index <= 2865) || (pixel_index >= 2895 && pixel_index <= 2960)) begin
            oled_data = PINK_HEX;
        end else if ((pixel_index >= 3705 && pixel_index <= 3707) || (pixel_index >= 3716 && pixel_index <= 3717) || (pixel_index >= 3801 && pixel_index <= 3803) || (pixel_index >= 3812 && pixel_index <= 3813) || (pixel_index >= 3897 && pixel_index <= 3899) || (pixel_index >= 3908 && pixel_index <= 3909) || (pixel_index >= 3958 && pixel_index <= 3959) || (pixel_index >= 3966 && pixel_index <= 3967) || (pixel_index >= 3972 && pixel_index <= 3977) || (pixel_index >= 3991 && pixel_index <= 3997) || (pixel_index >= 4004 && pixel_index <= 4005) || (pixel_index >= 4054 && pixel_index <= 4055) || (pixel_index >= 4062 && pixel_index <= 4063) || (pixel_index >= 4068 && pixel_index <= 4073) || (pixel_index >= 4087 && pixel_index <= 4088) || (pixel_index >= 4092 && pixel_index <= 4093) || (pixel_index >= 4100 && pixel_index <= 4101) || (pixel_index >= 4150 && pixel_index <= 4151) || (pixel_index >= 4158 && pixel_index <= 4159) || (pixel_index >= 4162 && pixel_index <= 4163) || (pixel_index >= 4183 && pixel_index <= 4184) || (pixel_index >= 4188 && pixel_index <= 4189) || (pixel_index >= 4196 && pixel_index <= 4197) || (pixel_index >= 4248 && pixel_index <= 4249) || (pixel_index >= 4252 && pixel_index <= 4253) || (pixel_index >= 4258 && pixel_index <= 4259) || (pixel_index >= 4278 && pixel_index <= 4280) || (pixel_index >= 4284 && pixel_index <= 4285) || (pixel_index >= 4292 && pixel_index <= 4293) || (pixel_index >= 4344 && pixel_index <= 4345) || (pixel_index >= 4348 && pixel_index <= 4349) || (pixel_index >= 4356 && pixel_index <= 4359) || (pixel_index >= 4374 && pixel_index <= 4382) || (pixel_index >= 4388 && pixel_index <= 4389) || (pixel_index >= 4440 && pixel_index <= 4441) || (pixel_index >= 4444 && pixel_index <= 4445) || (pixel_index >= 4452 && pixel_index <= 4455) || (pixel_index >= 4470 && pixel_index <= 4478) || (pixel_index >= 4484 && pixel_index <= 4485) || (pixel_index >= 4538 && pixel_index <= 4539) || (pixel_index >= 4552 && pixel_index <= 4553) || (pixel_index >= 4565 && pixel_index <= 4566) || (pixel_index >= 4574 && pixel_index <= 4575) || (pixel_index >= 4580 && pixel_index <= 4581) || (pixel_index >= 4634 && pixel_index <= 4635) || (pixel_index >= 4648 && pixel_index <= 4649) || (pixel_index >= 4661 && pixel_index <= 4662) || (pixel_index >= 4670 && pixel_index <= 4671) || (pixel_index >= 4676 && pixel_index <= 4677) || (pixel_index >= 4730 && pixel_index <= 4731) || (pixel_index >= 4738 && pixel_index <= 4743) || (pixel_index >= 4757 && pixel_index <= 4758) || (pixel_index >= 4766 && pixel_index <= 4767) || (pixel_index >= 4772 && pixel_index <= 4773) || (pixel_index >= 4826 && pixel_index <= 4827) || (pixel_index >= 4834 && pixel_index <= 4839) || (pixel_index >= 4853 && pixel_index <= 4854) || (pixel_index >= 4862 && pixel_index <= 4863) || (pixel_index >= 4868 && pixel_index <= 4869)) begin
            oled_data = BLUE_HEX;
        end else if ((pixel_index >= 1277 && pixel_index <= 1278) || (pixel_index >= 1313 && pixel_index <= 1314) || (pixel_index >= 1373 && pixel_index <= 1374) || (pixel_index >= 1409 && pixel_index <= 1410) || (pixel_index >= 1465 && pixel_index <= 1470) || (pixel_index >= 1501 && pixel_index <= 1506) || (pixel_index >= 1561 && pixel_index <= 1566) || (pixel_index >= 1578 && pixel_index <= 1579) || (pixel_index >= 1586 && pixel_index <= 1587) || (pixel_index >= 1597 && pixel_index <= 1602) || (pixel_index >= 1661 && pixel_index <= 1662) || (pixel_index >= 1674 && pixel_index <= 1675) || (pixel_index >= 1682 && pixel_index <= 1683) || (pixel_index >= 1697 && pixel_index <= 1698) || (pixel_index >= 1757 && pixel_index <= 1758) || (pixel_index >= 1772 && pixel_index <= 1773) || (pixel_index >= 1776 && pixel_index <= 1777) || (pixel_index >= 1793 && pixel_index <= 1794) || (pixel_index >= 1853 && pixel_index <= 1854) || (pixel_index >= 1868 && pixel_index <= 1869) || (pixel_index >= 1872 && pixel_index <= 1873) || (pixel_index >= 1889 && pixel_index <= 1890) || (pixel_index >= 1949 && pixel_index <= 1950) || (pixel_index >= 1964 && pixel_index <= 1965) || (pixel_index >= 1968 && pixel_index <= 1969) || (pixel_index >= 1985 && pixel_index <= 1986) || (pixel_index >= 2045 && pixel_index <= 2046) || (pixel_index >= 2060 && pixel_index <= 2061) || (pixel_index >= 2064 && pixel_index <= 2065) || (pixel_index >= 2081 && pixel_index <= 2082) || (pixel_index >= 2141 && pixel_index <= 2142) || (pixel_index >= 2158 && pixel_index <= 2159) || (pixel_index >= 2177 && pixel_index <= 2178) || (pixel_index >= 2237 && pixel_index <= 2238) || (pixel_index >= 2254 && pixel_index <= 2255) || (pixel_index >= 2273 && pixel_index <= 2274) || (pixel_index >= 2333 && pixel_index <= 2334) || (pixel_index >= 2350 && pixel_index <= 2351) || (pixel_index >= 2369 && pixel_index <= 2370) || (pixel_index >= 2429 && pixel_index <= 2430) || (pixel_index >= 2446 && pixel_index <= 2447) || (pixel_index >= 2465 && pixel_index <= 2466)) begin
            oled_data = WHITE_HEX;
        end else begin
            oled_data = BG_BLUE_HEX;
        end
    end    
endmodule

module display_mode_select_ai(
    input [12:0] pixel_index,
    output reg [15:0] oled_data
    );
    
    parameter PINK_HEX = 16'hF899;
    parameter BLUE_HEX = 16'h177F;
    parameter BG_BLUE_HEX = 16'h0006;
    parameter WHITE_HEX = 16'hFFFF;
    
    always @(*) begin
        if ((pixel_index >= 3087 && pixel_index <= 3152) || (pixel_index >= 3182 && pixel_index <= 3249) || (pixel_index >= 3277 && pixel_index <= 3346) || (pixel_index >= 3373 && pixel_index <= 3442) || (pixel_index >= 3469 && pixel_index <= 3538) || (pixel_index >= 3565 && pixel_index <= 3634) || (pixel_index >= 3661 && pixel_index <= 3704) || (pixel_index >= 3708 && pixel_index <= 3715) || (pixel_index >= 3718 && pixel_index <= 3730) || (pixel_index >= 3757 && pixel_index <= 3800) || (pixel_index >= 3804 && pixel_index <= 3811) || (pixel_index >= 3814 && pixel_index <= 3826) || (pixel_index >= 3853 && pixel_index <= 3896) || (pixel_index >= 3900 && pixel_index <= 3907) || (pixel_index >= 3910 && pixel_index <= 3922) || (pixel_index >= 3949 && pixel_index <= 3957) || (pixel_index >= 3960 && pixel_index <= 3965) || (pixel_index >= 3968 && pixel_index <= 3971) || (pixel_index >= 3978 && pixel_index <= 3992) || (pixel_index >= 3996 && pixel_index <= 4003) || (pixel_index >= 4006 && pixel_index <= 4018) || (pixel_index >= 4045 && pixel_index <= 4053) || (pixel_index >= 4056 && pixel_index <= 4061) || (pixel_index >= 4064 && pixel_index <= 4067) || (pixel_index >= 4074 && pixel_index <= 4086) || (pixel_index >= 4089 && pixel_index <= 4091) || (pixel_index >= 4094 && pixel_index <= 4099) || (pixel_index >= 4102 && pixel_index <= 4114) || (pixel_index >= 4141 && pixel_index <= 4151) || (pixel_index >= 4154 && pixel_index <= 4155) || (pixel_index >= 4158 && pixel_index <= 4161) || (pixel_index >= 4164 && pixel_index <= 4182) || (pixel_index >= 4185 && pixel_index <= 4187) || (pixel_index >= 4190 && pixel_index <= 4195) || (pixel_index >= 4198 && pixel_index <= 4210) || (pixel_index >= 4237 && pixel_index <= 4247) || (pixel_index >= 4250 && pixel_index <= 4251) || (pixel_index >= 4254 && pixel_index <= 4257) || (pixel_index >= 4260 && pixel_index <= 4278) || (pixel_index >= 4281 && pixel_index <= 4283) || (pixel_index >= 4286 && pixel_index <= 4291) || (pixel_index >= 4294 && pixel_index <= 4306) || (pixel_index >= 4333 && pixel_index <= 4343) || (pixel_index >= 4346 && pixel_index <= 4347) || (pixel_index >= 4350 && pixel_index <= 4355) || (pixel_index >= 4360 && pixel_index <= 4373) || (pixel_index >= 4383 && pixel_index <= 4387) || (pixel_index >= 4390 && pixel_index <= 4402) || (pixel_index >= 4429 && pixel_index <= 4439) || (pixel_index >= 4442 && pixel_index <= 4443) || (pixel_index >= 4446 && pixel_index <= 4451) || (pixel_index >= 4456 && pixel_index <= 4469) || (pixel_index >= 4479 && pixel_index <= 4483) || (pixel_index >= 4486 && pixel_index <= 4498) || (pixel_index >= 4525 && pixel_index <= 4537) || (pixel_index >= 4540 && pixel_index <= 4551) || (pixel_index >= 4554 && pixel_index <= 4564) || (pixel_index >= 4567 && pixel_index <= 4573) || (pixel_index >= 4576 && pixel_index <= 4579) || (pixel_index >= 4582 && pixel_index <= 4594) || (pixel_index >= 4621 && pixel_index <= 4633) || (pixel_index >= 4636 && pixel_index <= 4647) || (pixel_index >= 4650 && pixel_index <= 4660) || (pixel_index >= 4663 && pixel_index <= 4669) || (pixel_index >= 4672 && pixel_index <= 4675) || (pixel_index >= 4678 && pixel_index <= 4690) || (pixel_index >= 4717 && pixel_index <= 4729) || (pixel_index >= 4732 && pixel_index <= 4737) || (pixel_index >= 4744 && pixel_index <= 4756) || (pixel_index >= 4759 && pixel_index <= 4765) || (pixel_index >= 4768 && pixel_index <= 4771) || (pixel_index >= 4774 && pixel_index <= 4786) || (pixel_index >= 4813 && pixel_index <= 4825) || (pixel_index >= 4828 && pixel_index <= 4833) || (pixel_index >= 4840 && pixel_index <= 4852) || (pixel_index >= 4855 && pixel_index <= 4861) || (pixel_index >= 4864 && pixel_index <= 4867) || (pixel_index >= 4870 && pixel_index <= 4882) || (pixel_index >= 4909 && pixel_index <= 4978) || (pixel_index >= 5005 && pixel_index <= 5074) || (pixel_index >= 5101 && pixel_index <= 5170) || (pixel_index >= 5198 && pixel_index <= 5265) || (pixel_index >= 5295 && pixel_index <= 5360)) begin
            oled_data = PINK_HEX;
        end else if ((pixel_index >= 1277 && pixel_index <= 1278) || (pixel_index >= 1313 && pixel_index <= 1314) || (pixel_index >= 1373 && pixel_index <= 1374) || (pixel_index >= 1409 && pixel_index <= 1410) || (pixel_index >= 1465 && pixel_index <= 1470) || (pixel_index >= 1501 && pixel_index <= 1506) || (pixel_index >= 1561 && pixel_index <= 1566) || (pixel_index >= 1578 && pixel_index <= 1579) || (pixel_index >= 1586 && pixel_index <= 1587) || (pixel_index >= 1597 && pixel_index <= 1602) || (pixel_index >= 1661 && pixel_index <= 1662) || (pixel_index >= 1674 && pixel_index <= 1675) || (pixel_index >= 1682 && pixel_index <= 1683) || (pixel_index >= 1697 && pixel_index <= 1698) || (pixel_index >= 1757 && pixel_index <= 1758) || (pixel_index >= 1772 && pixel_index <= 1773) || (pixel_index >= 1776 && pixel_index <= 1777) || (pixel_index >= 1793 && pixel_index <= 1794) || (pixel_index >= 1853 && pixel_index <= 1854) || (pixel_index >= 1868 && pixel_index <= 1869) || (pixel_index >= 1872 && pixel_index <= 1873) || (pixel_index >= 1889 && pixel_index <= 1890) || (pixel_index >= 1949 && pixel_index <= 1950) || (pixel_index >= 1964 && pixel_index <= 1965) || (pixel_index >= 1968 && pixel_index <= 1969) || (pixel_index >= 1985 && pixel_index <= 1986) || (pixel_index >= 2045 && pixel_index <= 2046) || (pixel_index >= 2060 && pixel_index <= 2061) || (pixel_index >= 2064 && pixel_index <= 2065) || (pixel_index >= 2081 && pixel_index <= 2082) || (pixel_index >= 2141 && pixel_index <= 2142) || (pixel_index >= 2158 && pixel_index <= 2159) || (pixel_index >= 2177 && pixel_index <= 2178) || (pixel_index >= 2237 && pixel_index <= 2238) || (pixel_index >= 2254 && pixel_index <= 2255) || (pixel_index >= 2273 && pixel_index <= 2274) || (pixel_index >= 2333 && pixel_index <= 2334) || (pixel_index >= 2350 && pixel_index <= 2351) || (pixel_index >= 2369 && pixel_index <= 2370) || (pixel_index >= 2429 && pixel_index <= 2430) || (pixel_index >= 2446 && pixel_index <= 2447) || (pixel_index >= 2465 && pixel_index <= 2466)) begin
            oled_data = BLUE_HEX;
        end else if ((pixel_index >= 3705 && pixel_index <= 3707) || (pixel_index >= 3716 && pixel_index <= 3717) || (pixel_index >= 3801 && pixel_index <= 3803) || (pixel_index >= 3812 && pixel_index <= 3813) || (pixel_index >= 3897 && pixel_index <= 3899) || (pixel_index >= 3908 && pixel_index <= 3909) || (pixel_index >= 3958 && pixel_index <= 3959) || (pixel_index >= 3966 && pixel_index <= 3967) || (pixel_index >= 3972 && pixel_index <= 3977) || (pixel_index >= 3993 && pixel_index <= 3995) || (pixel_index >= 4004 && pixel_index <= 4005) || (pixel_index >= 4054 && pixel_index <= 4055) || (pixel_index >= 4062 && pixel_index <= 4063) || (pixel_index >= 4068 && pixel_index <= 4073) || (pixel_index >= 4087 && pixel_index <= 4088) || (pixel_index >= 4092 && pixel_index <= 4093) || (pixel_index >= 4100 && pixel_index <= 4101) || (pixel_index >= 4152 && pixel_index <= 4153) || (pixel_index >= 4156 && pixel_index <= 4157) || (pixel_index >= 4162 && pixel_index <= 4163) || (pixel_index >= 4183 && pixel_index <= 4184) || (pixel_index >= 4188 && pixel_index <= 4189) || (pixel_index >= 4196 && pixel_index <= 4197) || (pixel_index >= 4248 && pixel_index <= 4249) || (pixel_index >= 4252 && pixel_index <= 4253) || (pixel_index >= 4258 && pixel_index <= 4259) || (pixel_index >= 4279 && pixel_index <= 4280) || (pixel_index >= 4284 && pixel_index <= 4285) || (pixel_index >= 4292 && pixel_index <= 4293) || (pixel_index >= 4344 && pixel_index <= 4345) || (pixel_index >= 4348 && pixel_index <= 4349) || (pixel_index >= 4356 && pixel_index <= 4359) || (pixel_index >= 4374 && pixel_index <= 4382) || (pixel_index >= 4388 && pixel_index <= 4389) || (pixel_index >= 4440 && pixel_index <= 4441) || (pixel_index >= 4444 && pixel_index <= 4445) || (pixel_index >= 4452 && pixel_index <= 4455) || (pixel_index >= 4470 && pixel_index <= 4478) || (pixel_index >= 4484 && pixel_index <= 4485) || (pixel_index >= 4538 && pixel_index <= 4539) || (pixel_index >= 4552 && pixel_index <= 4553) || (pixel_index >= 4565 && pixel_index <= 4566) || (pixel_index >= 4574 && pixel_index <= 4575) || (pixel_index >= 4580 && pixel_index <= 4581) || (pixel_index >= 4634 && pixel_index <= 4635) || (pixel_index >= 4648 && pixel_index <= 4649) || (pixel_index >= 4661 && pixel_index <= 4662) || (pixel_index >= 4670 && pixel_index <= 4671) || (pixel_index >= 4676 && pixel_index <= 4677) || (pixel_index >= 4730 && pixel_index <= 4731) || (pixel_index >= 4738 && pixel_index <= 4743) || (pixel_index >= 4757 && pixel_index <= 4758) || (pixel_index >= 4766 && pixel_index <= 4767) || (pixel_index >= 4772 && pixel_index <= 4773) || (pixel_index >= 4826 && pixel_index <= 4827) || (pixel_index >= 4834 && pixel_index <= 4839) || (pixel_index >= 4853 && pixel_index <= 4854) || (pixel_index >= 4862 && pixel_index <= 4863) || (pixel_index >= 4868 && pixel_index <= 4869)) begin
            oled_data = WHITE_HEX;
        end else begin
            oled_data = BG_BLUE_HEX;
        end
    end    
endmodule  
