`timescale 1ns / 1ps

module vsbase_data(input [12:0] pixel_index, output reg [15:0] oled_data);
   
    always @ (*) begin
        if (((pixel_index >= 194) && (pixel_index <= 285)) || ((pixel_index >= 290) && (pixel_index <= 381)) || ((pixel_index >= 386) && (pixel_index <= 387)) || ((pixel_index >= 476) && (pixel_index <= 477)) || ((pixel_index >= 482) && (pixel_index <= 483)) || ((pixel_index >= 572) && (pixel_index <= 573)) || ((pixel_index >= 578) && (pixel_index <= 579)) || ((pixel_index >= 609) && (pixel_index <= 610)) || ((pixel_index >= 619) && (pixel_index <= 620)) || ((pixel_index >= 627) && (pixel_index <= 628)) || ((pixel_index >= 637) && (pixel_index <= 638)) || ((pixel_index >= 668) && (pixel_index <= 669)) || ((pixel_index >= 674) && (pixel_index <= 675)) || ((pixel_index >= 705) && (pixel_index <= 706)) || ((pixel_index >= 715) && (pixel_index <= 716)) || ((pixel_index >= 723) && (pixel_index <= 724)) || ((pixel_index >= 733) && (pixel_index <= 734)) || ((pixel_index >= 764) && (pixel_index <= 765)) || ((pixel_index >= 770) && (pixel_index <= 771)) || ((pixel_index >= 799) && (pixel_index <= 802)) || ((pixel_index >= 811) && (pixel_index <= 812)) || ((pixel_index >= 819) && (pixel_index <= 820)) || ((pixel_index >= 827) && (pixel_index <= 830)) || ((pixel_index >= 860) && (pixel_index <= 861)) || ((pixel_index >= 866) && (pixel_index <= 867)) || ((pixel_index >= 895) && (pixel_index <= 898)) || ((pixel_index >= 907) && (pixel_index <= 908)) || ((pixel_index >= 915) && (pixel_index <= 916)) || ((pixel_index >= 923) && (pixel_index <= 926)) || ((pixel_index >= 956) && (pixel_index <= 957)) || ((pixel_index >= 962) && (pixel_index <= 963)) || ((pixel_index >= 993) && (pixel_index <= 994)) || ((pixel_index >= 1005) && (pixel_index <= 1006)) || ((pixel_index >= 1009) && (pixel_index <= 1010)) || ((pixel_index >= 1021) && (pixel_index <= 1022)) || ((pixel_index >= 1052) && (pixel_index <= 1053)) || ((pixel_index >= 1058) && (pixel_index <= 1059)) || ((pixel_index >= 1089) && (pixel_index <= 1090)) || ((pixel_index >= 1101) && (pixel_index <= 1102)) || ((pixel_index >= 1105) && (pixel_index <= 1106)) || ((pixel_index >= 1117) && (pixel_index <= 1118)) || ((pixel_index >= 1148) && (pixel_index <= 1149)) || ((pixel_index >= 1154) && (pixel_index <= 1155)) || ((pixel_index >= 1185) && (pixel_index <= 1186)) || ((pixel_index >= 1197) && (pixel_index <= 1198)) || ((pixel_index >= 1201) && (pixel_index <= 1202)) || ((pixel_index >= 1213) && (pixel_index <= 1214)) || ((pixel_index >= 1244) && (pixel_index <= 1245)) || ((pixel_index >= 1250) && (pixel_index <= 1251)) || ((pixel_index >= 1281) && (pixel_index <= 1282)) || ((pixel_index >= 1293) && (pixel_index <= 1294)) || ((pixel_index >= 1297) && (pixel_index <= 1298)) || ((pixel_index >= 1309) && (pixel_index <= 1310)) || ((pixel_index >= 1340) && (pixel_index <= 1341)) || ((pixel_index >= 1346) && (pixel_index <= 1347)) || ((pixel_index >= 1375) && (pixel_index <= 1380)) || ((pixel_index >= 1391) && (pixel_index <= 1392)) || ((pixel_index >= 1403) && (pixel_index <= 1408)) || ((pixel_index >= 1436) && (pixel_index <= 1437)) || ((pixel_index >= 1442) && (pixel_index <= 1443)) || ((pixel_index >= 1471) && (pixel_index <= 1476)) || ((pixel_index >= 1487) && (pixel_index <= 1488)) || ((pixel_index >= 1499) && (pixel_index <= 1504)) || ((pixel_index >= 1532) && (pixel_index <= 1533)) || ((pixel_index >= 1538) && (pixel_index <= 1539)) || ((pixel_index >= 1628) && (pixel_index <= 1629)) || ((pixel_index >= 1634) && (pixel_index <= 1635)) || ((pixel_index >= 1724) && (pixel_index <= 1725)) || ((pixel_index >= 1730) && (pixel_index <= 1821)) || ((pixel_index >= 1826) && (pixel_index <= 1917)) || ((pixel_index >= 2221) && (pixel_index <= 2224)) || ((pixel_index >= 2229) && (pixel_index <= 2230)) || ((pixel_index >= 2235) && (pixel_index <= 2236)) || ((pixel_index >= 2239) && (pixel_index <= 2244)) || ((pixel_index >= 2249) && (pixel_index <= 2254)) || ((pixel_index >= 2259) && (pixel_index <= 2266)) || ((pixel_index >= 2269) && (pixel_index <= 2270)) || ((pixel_index >= 2275) && (pixel_index <= 2276)) || ((pixel_index >= 2279) && (pixel_index <= 2288)) || ((pixel_index >= 2317) && (pixel_index <= 2320)) || ((pixel_index >= 2325) && (pixel_index <= 2326)) || ((pixel_index >= 2331) && (pixel_index <= 2332)) || ((pixel_index >= 2335) && (pixel_index <= 2340)) || ((pixel_index >= 2345) && (pixel_index <= 2350)) || ((pixel_index >= 2355) && (pixel_index <= 2362)) || ((pixel_index >= 2365) && (pixel_index <= 2366)) || ((pixel_index >= 2371) && (pixel_index <= 2372)) || ((pixel_index >= 2375) && (pixel_index <= 2384)) || ((pixel_index >= 2387) && (pixel_index <= 2388)) || ((pixel_index >= 2411) && (pixel_index <= 2412)) || ((pixel_index >= 2417) && (pixel_index <= 2418)) || ((pixel_index >= 2421) && (pixel_index <= 2422)) || ((pixel_index >= 2427) && (pixel_index <= 2428)) || ((pixel_index >= 2431) && (pixel_index <= 2432)) || ((pixel_index >= 2437) && (pixel_index <= 2438)) || ((pixel_index >= 2441) && (pixel_index <= 2442)) || ((pixel_index >= 2447) && (pixel_index <= 2448)) || ((pixel_index >= 2451) && (pixel_index <= 2452)) || ((pixel_index >= 2461) && (pixel_index <= 2464)) || ((pixel_index >= 2467) && (pixel_index <= 2468)) || ((pixel_index >= 2475) && (pixel_index <= 2476)) || ((pixel_index >= 2483) && (pixel_index <= 2484)) || ((pixel_index >= 2507) && (pixel_index <= 2508)) || ((pixel_index >= 2513) && (pixel_index <= 2514)) || ((pixel_index >= 2517) && (pixel_index <= 2518)) || ((pixel_index >= 2523) && (pixel_index <= 2524)) || ((pixel_index >= 2527) && (pixel_index <= 2528)) || ((pixel_index >= 2533) && (pixel_index <= 2534)) || ((pixel_index >= 2537) && (pixel_index <= 2538)) || ((pixel_index >= 2543) && (pixel_index <= 2544)) || ((pixel_index >= 2547) && (pixel_index <= 2548)) || ((pixel_index >= 2557) && (pixel_index <= 2560)) || ((pixel_index >= 2563) && (pixel_index <= 2564)) || ((pixel_index >= 2571) && (pixel_index <= 2572)) || ((pixel_index >= 2603) && (pixel_index <= 2604)) || ((pixel_index >= 2613) && (pixel_index <= 2614)) || ((pixel_index >= 2619) && (pixel_index <= 2620)) || ((pixel_index >= 2623) && (pixel_index <= 2628)) || ((pixel_index >= 2633) && (pixel_index <= 2638)) || ((pixel_index >= 2643) && (pixel_index <= 2648)) || ((pixel_index >= 2653) && (pixel_index <= 2654)) || ((pixel_index >= 2657) && (pixel_index <= 2660)) || ((pixel_index >= 2667) && (pixel_index <= 2668)) || ((pixel_index >= 2699) && (pixel_index <= 2700)) || ((pixel_index >= 2709) && (pixel_index <= 2710)) || ((pixel_index >= 2715) && (pixel_index <= 2716)) || ((pixel_index >= 2719) && (pixel_index <= 2724)) || ((pixel_index >= 2729) && (pixel_index <= 2734)) || ((pixel_index >= 2739) && (pixel_index <= 2744)) || ((pixel_index >= 2749) && (pixel_index <= 2750)) || ((pixel_index >= 2753) && (pixel_index <= 2756)) || ((pixel_index >= 2763) && (pixel_index <= 2764)) || ((pixel_index >= 2795) && (pixel_index <= 2796)) || ((pixel_index >= 2801) && (pixel_index <= 2802)) || ((pixel_index >= 2805) && (pixel_index <= 2806)) || ((pixel_index >= 2811) && (pixel_index <= 2812)) || ((pixel_index >= 2815) && (pixel_index <= 2816)) || ((pixel_index >= 2819) && (pixel_index <= 2820)) || ((pixel_index >= 2825) && (pixel_index <= 2826)) || ((pixel_index >= 2829) && (pixel_index <= 2830)) || ((pixel_index >= 2835) && (pixel_index <= 2836)) || ((pixel_index >= 2845) && (pixel_index <= 2846)) || ((pixel_index >= 2851) && (pixel_index <= 2852)) || ((pixel_index >= 2859) && (pixel_index <= 2860)) || ((pixel_index >= 2891) && (pixel_index <= 2892)) || ((pixel_index >= 2897) && (pixel_index <= 2898)) || ((pixel_index >= 2901) && (pixel_index <= 2902)) || ((pixel_index >= 2907) && (pixel_index <= 2908)) || ((pixel_index >= 2911) && (pixel_index <= 2912)) || ((pixel_index >= 2915) && (pixel_index <= 2916)) || ((pixel_index >= 2921) && (pixel_index <= 2922)) || ((pixel_index >= 2925) && (pixel_index <= 2926)) || ((pixel_index >= 2931) && (pixel_index <= 2932)) || ((pixel_index >= 2941) && (pixel_index <= 2942)) || ((pixel_index >= 2947) && (pixel_index <= 2948)) || ((pixel_index >= 2955) && (pixel_index <= 2956)) || ((pixel_index >= 2963) && (pixel_index <= 2964)) || ((pixel_index >= 2989) && (pixel_index <= 2992)) || ((pixel_index >= 2999) && (pixel_index <= 3002)) || ((pixel_index >= 3007) && (pixel_index <= 3008)) || ((pixel_index >= 3013) && (pixel_index <= 3014)) || ((pixel_index >= 3017) && (pixel_index <= 3018)) || ((pixel_index >= 3023) && (pixel_index <= 3024)) || ((pixel_index >= 3027) && (pixel_index <= 3034)) || ((pixel_index >= 3037) && (pixel_index <= 3038)) || ((pixel_index >= 3043) && (pixel_index <= 3044)) || ((pixel_index >= 3051) && (pixel_index <= 3052)) || ((pixel_index >= 3059) && (pixel_index <= 3060)) || ((pixel_index >= 3085) && (pixel_index <= 3088)) || ((pixel_index >= 3095) && (pixel_index <= 3098)) || ((pixel_index >= 3103) && (pixel_index <= 3104)) || ((pixel_index >= 3109) && (pixel_index <= 3110)) || ((pixel_index >= 3113) && (pixel_index <= 3114)) || ((pixel_index >= 3119) && (pixel_index <= 3120)) || ((pixel_index >= 3123) && (pixel_index <= 3130)) || ((pixel_index >= 3133) && (pixel_index <= 3134)) || ((pixel_index >= 3139) && (pixel_index <= 3140)) || (pixel_index >= 3147) && (pixel_index <= 3148)) oled_data = 16'b1111111111111111;
        else if (pixel_index >= 3264) oled_data = 0;
        else oled_data = 16'b0000000001000100;
    end

endmodule

module vsturn_data(input sw, input [12:0] pixel_index, output reg [15:0] oled_data);
   
    always @ (*) begin
        if (pixel_index <= 3263) oled_data = 0;
        if (sw == 0) begin // cross
            if (pixel_index == 3493 || pixel_index == 3513 || pixel_index == 3611 || pixel_index == 3689 || pixel_index == 3799 || pixel_index == 3893 || pixel_index == 3988 || pixel_index == 4086 || pixel_index == 4088 || pixel_index == 4277 || pixel_index == 4364 || pixel_index == 4368 || pixel_index == 4370 || pixel_index == 4560 || pixel_index == 4654 || pixel_index == 4844 || pixel_index == 4852 || pixel_index == 4945 || pixel_index == 4949 || pixel_index == 5034 || pixel_index == 5036 || pixel_index == 5228 || pixel_index == 5235 || pixel_index == 5623 || pixel_index == 5722 || pixel_index == 5724 || pixel_index == 5799 || pixel_index == 3494 || pixel_index == 3514 || pixel_index == 3589 || ((pixel_index >= 3609) && (pixel_index <= 3610)) || pixel_index == 3612 || pixel_index == 3684 || ((pixel_index >= 3687) && (pixel_index <= 3688)) || pixel_index == 3703 || pixel_index == 3707 || pixel_index == 3781 || pixel_index == 3785 || pixel_index == 3798 || pixel_index == 3802 || pixel_index == 3804 || pixel_index == 3879 || pixel_index == 3883 || pixel_index == 3894 || pixel_index == 3896 || pixel_index == 3899 || pixel_index == 3974 || pixel_index == 3976 || pixel_index == 3978 || pixel_index == 3989 || pixel_index == 3991 || pixel_index == 3993 || pixel_index == 4075 || ((pixel_index >= 4084) && (pixel_index <= 4085)) || pixel_index == 4087 || ((pixel_index >= 4168) && (pixel_index <= 4169)) || ((pixel_index >= 4173) && (pixel_index <= 4174)) || pixel_index == 4178 || pixel_index == 4181 || pixel_index == 4184 || pixel_index == 4268 || pixel_index == 4274 || pixel_index == 4276 || pixel_index == 4278 || pixel_index == 4363 || pixel_index == 4365 || pixel_index == 4367 || pixel_index == 4369 || pixel_index == 4371 || pixel_index == 4373 || pixel_index == 4460 || ((pixel_index >= 4464) && (pixel_index <= 4465)) || pixel_index == 4467 || ((pixel_index >= 4556) && (pixel_index <= 4557)) || pixel_index == 4559 || pixel_index == 4561 || pixel_index == 4653 || pixel_index == 4655 || pixel_index == 4657 || pixel_index == 4659 || pixel_index == 4749 || pixel_index == 4751 || pixel_index == 4756 || pixel_index == 4843 || pixel_index == 4845 || pixel_index == 4848 || ((pixel_index >= 4850) && (pixel_index <= 4851)) || pixel_index == 4853 || pixel_index == 4938 || pixel_index == 4940 || pixel_index == 4944 || pixel_index == 4946 || pixel_index == 4948 || pixel_index == 4950 || pixel_index == 5033 || pixel_index == 5035 || pixel_index == 5037 || pixel_index == 5041 || pixel_index == 5045 || pixel_index == 5047 || pixel_index == 5130 || ((pixel_index >= 5139) && (pixel_index <= 5140)) || pixel_index == 5144 || ((pixel_index >= 5223) && (pixel_index <= 5224)) || pixel_index == 5227 || pixel_index == 5229 || pixel_index == 5236 || pixel_index == 5241 || pixel_index == 5318 || pixel_index == 5320 || pixel_index == 5322 || pixel_index == 5324 || pixel_index == 5332 || pixel_index == 5335 || pixel_index == 5413 || pixel_index == 5429 || pixel_index == 5433 || pixel_index == 5435 || pixel_index == 5511 || ((pixel_index >= 5513) && (pixel_index <= 5514)) || ((pixel_index >= 5527) && (pixel_index <= 5528)) || pixel_index == 5530 || pixel_index == 5604 || pixel_index == 5606 || pixel_index == 5624 || ((pixel_index >= 5626) && (pixel_index <= 5627)) || ((pixel_index >= 5703) && (pixel_index <= 5704)) || ((pixel_index >= 5720) && (pixel_index <= 5721)) || pixel_index == 5723 || ((pixel_index >= 5797) && (pixel_index <= 5798)) || pixel_index == 5818 || pixel_index == 3495 || pixel_index == 3515 || pixel_index == 3588 || pixel_index == 3590 || pixel_index == 3592 || pixel_index == 3608 || pixel_index == 3686 || pixel_index == 3704 || pixel_index == 3706 || pixel_index == 3708 || pixel_index == 3780 || pixel_index == 3782 || pixel_index == 3784 || pixel_index == 3786 || pixel_index == 3801 || pixel_index == 3880 || pixel_index == 3882 || pixel_index == 3895 || pixel_index == 3898 || pixel_index == 3975 || pixel_index == 3980 || pixel_index == 3990 || pixel_index == 3992 || pixel_index == 3994 || pixel_index == 4072 || pixel_index == 4074 || pixel_index == 4076 || pixel_index == 4083 || pixel_index == 4170 || pixel_index == 4172 || pixel_index == 4180 || pixel_index == 4182 || pixel_index == 4266 || pixel_index == 4269 || pixel_index == 4271 || pixel_index == 4273 || pixel_index == 4275 || pixel_index == 4279 || pixel_index == 4362 || pixel_index == 4366 || pixel_index == 4372 || pixel_index == 4374 || pixel_index == 4459 || pixel_index == 4461 || pixel_index == 4463 || pixel_index == 4466 || pixel_index == 4469 || pixel_index == 4558 || pixel_index == 4564 || pixel_index == 4656 || pixel_index == 4658 || pixel_index == 4748 || pixel_index == 4750 || pixel_index == 4753 || pixel_index == 4755 || pixel_index == 4847 || pixel_index == 4849 || pixel_index == 4939 || pixel_index == 4941 || pixel_index == 4943 || pixel_index == 4947 || pixel_index == 5038 || pixel_index == 5042 || pixel_index == 5044 || pixel_index == 5046 || pixel_index == 5131 || pixel_index == 5133 || pixel_index == 5138 || pixel_index == 5141 || pixel_index == 5143 || pixel_index == 5225 || pixel_index == 5237 || pixel_index == 5239 || pixel_index == 5319 || pixel_index == 5321 || pixel_index == 5323 || pixel_index == 5334 || pixel_index == 5336 || pixel_index == 5338 || pixel_index == 5414 || pixel_index == 5418 || pixel_index == 5430 || pixel_index == 5432 || pixel_index == 5434 || pixel_index == 5508 || pixel_index == 5510 || pixel_index == 5512 || pixel_index == 5526 || pixel_index == 5531 || pixel_index == 5605 || pixel_index == 5607 || pixel_index == 5609 || pixel_index == 5625 || pixel_index == 5628 || pixel_index == 5700 || pixel_index == 5817 || pixel_index == 3591 || pixel_index == 3685 || pixel_index == 3705 || pixel_index == 3783 || pixel_index == 3877 || pixel_index == 3881 || pixel_index == 3897 || pixel_index == 3979 || pixel_index == 4071 || pixel_index == 4073 || pixel_index == 4077 || pixel_index == 4171 || pixel_index == 4179 || pixel_index == 4265 || pixel_index == 4270 || pixel_index == 4563 || pixel_index == 4754 || pixel_index == 4846 || pixel_index == 5039 || pixel_index == 5128 || pixel_index == 5134 || pixel_index == 5142 || pixel_index == 5226 || pixel_index == 5240 || pixel_index == 5333 || pixel_index == 5337 || pixel_index == 5415 || pixel_index == 5417 || pixel_index == 5431 || pixel_index == 5509 || pixel_index == 5532 || pixel_index == 5608 || pixel_index == 5701 || pixel_index == 3800 || pixel_index == 4089 || pixel_index == 4183 || pixel_index == 4267 || pixel_index == 4942 || pixel_index == 5132 || pixel_index == 5238 || pixel_index == 5419 || pixel_index == 3803 || pixel_index == 5529 || pixel_index == 3878 || pixel_index == 3977 || pixel_index == 4562 || pixel_index == 5129 || pixel_index == 5416 || pixel_index == 5702 || pixel_index == 5819 || pixel_index == 4462 || pixel_index == 4468 || pixel_index == 4752 || pixel_index == 5043) oled_data = 16'b0001011101111111;
            else oled_data = 16'b0000000001000100;
        end
        if (sw == 1) begin // circle
            if (((pixel_index >= 3403) && (pixel_index <= 3404)) || ((pixel_index >= 3406) && (pixel_index <= 3407)) || pixel_index == 3409 || pixel_index == 3412 || pixel_index == 3501 || pixel_index == 3504 || pixel_index == 3506 || pixel_index == 3510 || pixel_index == 3593 || ((pixel_index >= 3595) && (pixel_index <= 3596)) || pixel_index == 3598 || pixel_index == 3600 || ((pixel_index >= 3602) && (pixel_index <= 3603)) || pixel_index == 3687 || ((pixel_index >= 3692) && (pixel_index <= 3693)) || pixel_index == 3697 || ((pixel_index >= 3701) && (pixel_index <= 3702)) || pixel_index == 3704 || pixel_index == 3783 || ((pixel_index >= 3785) && (pixel_index <= 3786)) || ((pixel_index >= 3795) && (pixel_index <= 3796)) || pixel_index == 3798 || pixel_index == 3878 || pixel_index == 3880 || pixel_index == 3882 || pixel_index == 3893 || pixel_index == 3895 || ((pixel_index >= 3897) && (pixel_index <= 3898)) || pixel_index == 3973 || pixel_index == 3975 || pixel_index == 3977 || pixel_index == 3991 || pixel_index == 4070 || pixel_index == 4073 || pixel_index == 4086 || pixel_index == 4088 || ((pixel_index >= 4090) && (pixel_index <= 4091)) || ((pixel_index >= 4163) && (pixel_index <= 4164)) || pixel_index == 4166 || pixel_index == 4168 || pixel_index == 4260 || ((pixel_index >= 4262) && (pixel_index <= 4263)) || ((pixel_index >= 4280) && (pixel_index <= 4281)) || pixel_index == 4283 || pixel_index == 4355 || pixel_index == 4357 || pixel_index == 4359 || pixel_index == 4376 || pixel_index == 4378 || pixel_index == 4380 || pixel_index == 4452 || ((pixel_index >= 4474) && (pixel_index <= 4475)) || pixel_index == 4547 || pixel_index == 4549 || pixel_index == 4572 || pixel_index == 4643 || pixel_index == 4646 || ((pixel_index >= 4665) && (pixel_index <= 4666)) || pixel_index == 4668 || pixel_index == 4739 || pixel_index == 4741 || pixel_index == 4762 || pixel_index == 4764 || pixel_index == 4836 || pixel_index == 4838 || pixel_index == 4859 || pixel_index == 4932 || pixel_index == 4934 || ((pixel_index >= 4952) && (pixel_index <= 4953)) || pixel_index == 4956 || ((pixel_index >= 5028) && (pixel_index <= 5029)) || pixel_index == 5031 || pixel_index == 5047 || ((pixel_index >= 5049) && (pixel_index <= 5050)) || pixel_index == 5052 || pixel_index == 5124 || pixel_index == 5126 || pixel_index == 5143 || pixel_index == 5145 || pixel_index == 5147 || pixel_index == 5220 || pixel_index == 5222 || pixel_index == 5225 || pixel_index == 5237 || pixel_index == 5239 || pixel_index == 5241 || pixel_index == 5243 || ((pixel_index >= 5319) && (pixel_index <= 5320)) || pixel_index == 5322 || pixel_index == 5335 || pixel_index == 5337 || pixel_index == 5414 || pixel_index == 5416 || pixel_index == 5418 || pixel_index == 5427 || pixel_index == 5429 || pixel_index == 5431 || pixel_index == 5510 || pixel_index == 5512 || pixel_index == 5514 || pixel_index == 5516 || pixel_index == 5518 || ((pixel_index >= 5520) && (pixel_index <= 5521)) || pixel_index == 5523 || pixel_index == 5526 || pixel_index == 5528 || pixel_index == 5609 || pixel_index == 5612 || ((pixel_index >= 5614) && (pixel_index <= 5615)) || pixel_index == 5619 || pixel_index == 5622 || pixel_index == 5706 || ((pixel_index >= 5708) && (pixel_index <= 5709)) || pixel_index == 5713 || pixel_index == 5715 || pixel_index == 5717 || pixel_index == 5803 || pixel_index == 5805 || pixel_index == 5807 || (pixel_index >= 5809) && (pixel_index <= 5810) || pixel_index == 3405 || pixel_index == 3597 || pixel_index == 3601 || pixel_index == 3686 || pixel_index == 3797 || pixel_index == 3879 || pixel_index == 3881 || pixel_index == 4167 || pixel_index == 4259 || pixel_index == 4261 || pixel_index == 4377 || pixel_index == 4379 || pixel_index == 4451 || pixel_index == 4763 || pixel_index == 4933 || pixel_index == 5027 || pixel_index == 5048 || pixel_index == 5125 || pixel_index == 5146 || pixel_index == 5240 || pixel_index == 5415 || pixel_index == 5417 || pixel_index == 5519 || pixel_index == 5613 || pixel_index == 5623 || pixel_index == 5714 || pixel_index == 5804 || pixel_index == 3408 || pixel_index == 3411 || pixel_index == 3498 || pixel_index == 3500 || pixel_index == 3502 || pixel_index == 3505 || pixel_index == 3507 || pixel_index == 3509 || pixel_index == 3592 || pixel_index == 3594 || pixel_index == 3599 || pixel_index == 3604 || pixel_index == 3606 || pixel_index == 3689 || pixel_index == 3691 || pixel_index == 3694 || pixel_index == 3696 || pixel_index == 3698 || pixel_index == 3700 || pixel_index == 3703 || pixel_index == 3782 || pixel_index == 3784 || pixel_index == 3787 || pixel_index == 3789 || pixel_index == 3794 || pixel_index == 3799 || pixel_index == 3801 || pixel_index == 3883 || pixel_index == 3892 || pixel_index == 3894 || pixel_index == 3896 || pixel_index == 3972 || pixel_index == 3974 || pixel_index == 3976 || pixel_index == 3978 || pixel_index == 3989 || pixel_index == 3993 || pixel_index == 3995 || pixel_index == 4068 || pixel_index == 4071 || pixel_index == 4087 || pixel_index == 4089 || pixel_index == 4165 || pixel_index == 4184 || pixel_index == 4186 || pixel_index == 4188 || pixel_index == 4282 || pixel_index == 4284 || pixel_index == 4356 || pixel_index == 4358 || pixel_index == 4454 || pixel_index == 4473 || pixel_index == 4476 || pixel_index == 4548 || pixel_index == 4550 || pixel_index == 4570 || pixel_index == 4645 || pixel_index == 4667 || pixel_index == 4740 || pixel_index == 4761 || pixel_index == 4837 || pixel_index == 4839 || pixel_index == 4856 || pixel_index == 4858 || pixel_index == 4860 || pixel_index == 4931 || pixel_index == 4954 || pixel_index == 5030 || pixel_index == 5032 || pixel_index == 5051 || pixel_index == 5127 || pixel_index == 5129 || pixel_index == 5144 || pixel_index == 5221 || pixel_index == 5224 || pixel_index == 5238 || pixel_index == 5242 || pixel_index == 5318 || pixel_index == 5321 || pixel_index == 5323 || pixel_index == 5333 || pixel_index == 5336 || pixel_index == 5420 || pixel_index == 5428 || pixel_index == 5430 || pixel_index == 5433 || pixel_index == 5511 || pixel_index == 5513 || pixel_index == 5515 || pixel_index == 5517 || pixel_index == 5522 || pixel_index == 5525 || pixel_index == 5527 || pixel_index == 5529 || pixel_index == 5610 || pixel_index == 5616 || pixel_index == 5618 || pixel_index == 5620 || pixel_index == 5705 || pixel_index == 5707 || pixel_index == 5710 || pixel_index == 5712 || pixel_index == 5716 || pixel_index == 5718 || pixel_index == 5806 || pixel_index == 5808 || pixel_index == 5811 || pixel_index == 3410 || pixel_index == 3497 || pixel_index == 3499 || pixel_index == 3503 || pixel_index == 3508 || pixel_index == 3605 || pixel_index == 3607 || pixel_index == 3688 || pixel_index == 3690 || pixel_index == 3695 || pixel_index == 3699 || pixel_index == 3705 || pixel_index == 3788 || pixel_index == 3800 || pixel_index == 3877 || pixel_index == 3990 || pixel_index == 3992 || pixel_index == 3994 || pixel_index == 4069 || pixel_index == 4072 || pixel_index == 4183 || pixel_index == 4185 || pixel_index == 4187 || pixel_index == 4453 || pixel_index == 4569 || pixel_index == 4571 || pixel_index == 4644 || pixel_index == 4742 || pixel_index == 4835 || pixel_index == 4857 || pixel_index == 4935 || pixel_index == 4955 || pixel_index == 5128 || pixel_index == 5142 || pixel_index == 5223 || pixel_index == 5226 || pixel_index == 5317 || pixel_index == 5332 || pixel_index == 5334 || pixel_index == 5338 || pixel_index == 5419 || pixel_index == 5421 || pixel_index == 5426 || pixel_index == 5432 || pixel_index == 5524 || pixel_index == 5608 || pixel_index == 5611 || pixel_index == 5617 || pixel_index == 5621 || pixel_index == 5711 || pixel_index == 5812) oled_data = 16'b1111100001011010;
            else oled_data = 16'b0000000001000100;
        end
    end

endmodule