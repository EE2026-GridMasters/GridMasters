`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05/18/2024 05:51:42 PM
// Design Name: 
// Module Name: frame_data
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module airesult_data(input [1:0] result, input [12:0] pixel_index, output reg [15:0] oled_data);

    always @ (*) begin
        if (result == 2'b00) oled_data = 0;
        else if (result == 2'b01) begin // player win
            if (((pixel_index >= 194) && (pixel_index <= 285)) || ((pixel_index >= 290) && (pixel_index <= 381)) || ((pixel_index >= 386) && (pixel_index <= 387)) || ((pixel_index >= 476) && (pixel_index <= 477)) || ((pixel_index >= 482) && (pixel_index <= 483)) || ((pixel_index >= 572) && (pixel_index <= 573)) || ((pixel_index >= 578) && (pixel_index <= 579)) || ((pixel_index >= 592) && (pixel_index <= 593)) || ((pixel_index >= 600) && (pixel_index <= 601)) || ((pixel_index >= 606) && (pixel_index <= 609)) || ((pixel_index >= 614) && (pixel_index <= 615)) || ((pixel_index >= 620) && (pixel_index <= 621)) || ((pixel_index >= 668) && (pixel_index <= 669)) || ((pixel_index >= 674) && (pixel_index <= 675)) || ((pixel_index >= 688) && (pixel_index <= 689)) || ((pixel_index >= 696) && (pixel_index <= 697)) || ((pixel_index >= 702) && (pixel_index <= 705)) || ((pixel_index >= 710) && (pixel_index <= 711)) || ((pixel_index >= 716) && (pixel_index <= 717)) || ((pixel_index >= 764) && (pixel_index <= 765)) || ((pixel_index >= 770) && (pixel_index <= 771)) || ((pixel_index >= 784) && (pixel_index <= 785)) || ((pixel_index >= 792) && (pixel_index <= 793)) || ((pixel_index >= 796) && (pixel_index <= 797)) || ((pixel_index >= 802) && (pixel_index <= 803)) || ((pixel_index >= 806) && (pixel_index <= 807)) || ((pixel_index >= 812) && (pixel_index <= 813)) || ((pixel_index >= 860) && (pixel_index <= 861)) || ((pixel_index >= 866) && (pixel_index <= 867)) || ((pixel_index >= 880) && (pixel_index <= 881)) || ((pixel_index >= 888) && (pixel_index <= 889)) || ((pixel_index >= 892) && (pixel_index <= 893)) || ((pixel_index >= 898) && (pixel_index <= 899)) || ((pixel_index >= 902) && (pixel_index <= 903)) || ((pixel_index >= 908) && (pixel_index <= 909)) || ((pixel_index >= 956) && (pixel_index <= 957)) || ((pixel_index >= 962) && (pixel_index <= 963)) || ((pixel_index >= 978) && (pixel_index <= 983)) || ((pixel_index >= 988) && (pixel_index <= 989)) || ((pixel_index >= 994) && (pixel_index <= 995)) || ((pixel_index >= 998) && (pixel_index <= 999)) || ((pixel_index >= 1004) && (pixel_index <= 1005)) || ((pixel_index >= 1052) && (pixel_index <= 1053)) || ((pixel_index >= 1058) && (pixel_index <= 1059)) || ((pixel_index >= 1074) && (pixel_index <= 1079)) || ((pixel_index >= 1084) && (pixel_index <= 1085)) || ((pixel_index >= 1090) && (pixel_index <= 1091)) || ((pixel_index >= 1094) && (pixel_index <= 1095)) || ((pixel_index >= 1100) && (pixel_index <= 1101)) || ((pixel_index >= 1148) && (pixel_index <= 1149)) || ((pixel_index >= 1154) && (pixel_index <= 1155)) || ((pixel_index >= 1172) && (pixel_index <= 1173)) || ((pixel_index >= 1180) && (pixel_index <= 1181)) || ((pixel_index >= 1186) && (pixel_index <= 1187)) || ((pixel_index >= 1190) && (pixel_index <= 1191)) || ((pixel_index >= 1196) && (pixel_index <= 1197)) || ((pixel_index >= 1244) && (pixel_index <= 1245)) || ((pixel_index >= 1250) && (pixel_index <= 1251)) || ((pixel_index >= 1268) && (pixel_index <= 1269)) || ((pixel_index >= 1276) && (pixel_index <= 1277)) || ((pixel_index >= 1282) && (pixel_index <= 1283)) || ((pixel_index >= 1286) && (pixel_index <= 1287)) || ((pixel_index >= 1292) && (pixel_index <= 1293)) || ((pixel_index >= 1340) && (pixel_index <= 1341)) || ((pixel_index >= 1346) && (pixel_index <= 1347)) || ((pixel_index >= 1364) && (pixel_index <= 1365)) || ((pixel_index >= 1374) && (pixel_index <= 1377)) || ((pixel_index >= 1384) && (pixel_index <= 1387)) || ((pixel_index >= 1436) && (pixel_index <= 1437)) || ((pixel_index >= 1442) && (pixel_index <= 1443)) || ((pixel_index >= 1460) && (pixel_index <= 1461)) || ((pixel_index >= 1470) && (pixel_index <= 1473)) || ((pixel_index >= 1480) && (pixel_index <= 1483)) || ((pixel_index >= 1532) && (pixel_index <= 1533)) || ((pixel_index >= 1538) && (pixel_index <= 1539)) || ((pixel_index >= 1628) && (pixel_index <= 1629)) || ((pixel_index >= 1634) && (pixel_index <= 1635)) || ((pixel_index >= 1724) && (pixel_index <= 1725)) || ((pixel_index >= 1730) && (pixel_index <= 1821)) || ((pixel_index >= 1826) && (pixel_index <= 1917)) || ((pixel_index >= 3700) && (pixel_index <= 3701)) || ((pixel_index >= 3706) && (pixel_index <= 3707)) || ((pixel_index >= 3710) && (pixel_index <= 3717)) || ((pixel_index >= 3720) && (pixel_index <= 3721)) || ((pixel_index >= 3726) && (pixel_index <= 3727)) || ((pixel_index >= 3730) && (pixel_index <= 3739)) || ((pixel_index >= 3796) && (pixel_index <= 3797)) || ((pixel_index >= 3802) && (pixel_index <= 3803)) || ((pixel_index >= 3806) && (pixel_index <= 3813)) || ((pixel_index >= 3816) && (pixel_index <= 3817)) || ((pixel_index >= 3822) && (pixel_index <= 3823)) || ((pixel_index >= 3826) && (pixel_index <= 3835)) || ((pixel_index >= 3892) && (pixel_index <= 3895)) || ((pixel_index >= 3898) && (pixel_index <= 3899)) || ((pixel_index >= 3902) && (pixel_index <= 3903)) || ((pixel_index >= 3912) && (pixel_index <= 3913)) || ((pixel_index >= 3918) && (pixel_index <= 3919)) || ((pixel_index >= 3926) && (pixel_index <= 3927)) || ((pixel_index >= 3988) && (pixel_index <= 3991)) || ((pixel_index >= 3994) && (pixel_index <= 3995)) || ((pixel_index >= 3998) && (pixel_index <= 3999)) || ((pixel_index >= 4008) && (pixel_index <= 4009)) || ((pixel_index >= 4014) && (pixel_index <= 4015)) || ((pixel_index >= 4022) && (pixel_index <= 4023)) || ((pixel_index >= 4084) && (pixel_index <= 4085)) || ((pixel_index >= 4088) && (pixel_index <= 4091)) || ((pixel_index >= 4094) && (pixel_index <= 4099)) || ((pixel_index >= 4106) && (pixel_index <= 4109)) || ((pixel_index >= 4118) && (pixel_index <= 4119)) || ((pixel_index >= 4180) && (pixel_index <= 4181)) || ((pixel_index >= 4184) && (pixel_index <= 4187)) || ((pixel_index >= 4190) && (pixel_index <= 4195)) || ((pixel_index >= 4202) && (pixel_index <= 4205)) || ((pixel_index >= 4214) && (pixel_index <= 4215)) || ((pixel_index >= 4276) && (pixel_index <= 4277)) || ((pixel_index >= 4282) && (pixel_index <= 4283)) || ((pixel_index >= 4286) && (pixel_index <= 4287)) || ((pixel_index >= 4296) && (pixel_index <= 4297)) || ((pixel_index >= 4302) && (pixel_index <= 4303)) || ((pixel_index >= 4310) && (pixel_index <= 4311)) || ((pixel_index >= 4372) && (pixel_index <= 4373)) || ((pixel_index >= 4378) && (pixel_index <= 4379)) || ((pixel_index >= 4382) && (pixel_index <= 4383)) || ((pixel_index >= 4392) && (pixel_index <= 4393)) || ((pixel_index >= 4398) && (pixel_index <= 4399)) || ((pixel_index >= 4406) && (pixel_index <= 4407)) || ((pixel_index >= 4468) && (pixel_index <= 4469)) || ((pixel_index >= 4474) && (pixel_index <= 4475)) || ((pixel_index >= 4478) && (pixel_index <= 4485)) || ((pixel_index >= 4488) && (pixel_index <= 4489)) || ((pixel_index >= 4494) && (pixel_index <= 4495)) || ((pixel_index >= 4502) && (pixel_index <= 4503)) || ((pixel_index >= 4564) && (pixel_index <= 4565)) || ((pixel_index >= 4570) && (pixel_index <= 4571)) || ((pixel_index >= 4574) && (pixel_index <= 4581)) || ((pixel_index >= 4584) && (pixel_index <= 4585)) || ((pixel_index >= 4590) && (pixel_index <= 4591)) || ((pixel_index >= 4598) && (pixel_index <= 4599)) || ((pixel_index >= 4831) && (pixel_index <= 4832)) || ((pixel_index >= 4842) && (pixel_index <= 4843)) || ((pixel_index >= 4852) && (pixel_index <= 4859)) || ((pixel_index >= 4862) && (pixel_index <= 4863)) || ((pixel_index >= 4870) && (pixel_index <= 4871)) || ((pixel_index >= 4874) && (pixel_index <= 4881)) || ((pixel_index >= 4884) && (pixel_index <= 4885)) || ((pixel_index >= 4927) && (pixel_index <= 4929)) || ((pixel_index >= 4938) && (pixel_index <= 4939)) || ((pixel_index >= 4948) && (pixel_index <= 4955)) || ((pixel_index >= 4958) && (pixel_index <= 4959)) || ((pixel_index >= 4966) && (pixel_index <= 4967)) || ((pixel_index >= 4970) && (pixel_index <= 4977)) || ((pixel_index >= 4980) && (pixel_index <= 4981)) || ((pixel_index >= 5024) && (pixel_index <= 5026)) || ((pixel_index >= 5034) && (pixel_index <= 5035)) || ((pixel_index >= 5044) && (pixel_index <= 5045)) || ((pixel_index >= 5054) && (pixel_index <= 5055)) || ((pixel_index >= 5062) && (pixel_index <= 5063)) || ((pixel_index >= 5066) && (pixel_index <= 5067)) || ((pixel_index >= 5076) && (pixel_index <= 5077)) || ((pixel_index >= 5121) && (pixel_index <= 5123)) || ((pixel_index >= 5130) && (pixel_index <= 5131)) || ((pixel_index >= 5140) && (pixel_index <= 5141)) || ((pixel_index >= 5150) && (pixel_index <= 5151)) || ((pixel_index >= 5158) && (pixel_index <= 5159)) || ((pixel_index >= 5162) && (pixel_index <= 5163)) || ((pixel_index >= 5172) && (pixel_index <= 5173)) || ((pixel_index >= 5205) && (pixel_index <= 5220)) || ((pixel_index >= 5226) && (pixel_index <= 5227)) || ((pixel_index >= 5236) && (pixel_index <= 5241)) || ((pixel_index >= 5248) && (pixel_index <= 5249)) || ((pixel_index >= 5252) && (pixel_index <= 5253)) || ((pixel_index >= 5258) && (pixel_index <= 5263)) || ((pixel_index >= 5268) && (pixel_index <= 5269)) || ((pixel_index >= 5301) && (pixel_index <= 5316)) || ((pixel_index >= 5322) && (pixel_index <= 5323)) || ((pixel_index >= 5332) && (pixel_index <= 5337)) || ((pixel_index >= 5344) && (pixel_index <= 5345)) || ((pixel_index >= 5348) && (pixel_index <= 5349)) || ((pixel_index >= 5354) && (pixel_index <= 5359)) || ((pixel_index >= 5364) && (pixel_index <= 5365)) || ((pixel_index >= 5409) && (pixel_index <= 5411)) || ((pixel_index >= 5418) && (pixel_index <= 5419)) || ((pixel_index >= 5428) && (pixel_index <= 5429)) || ((pixel_index >= 5440) && (pixel_index <= 5441)) || ((pixel_index >= 5444) && (pixel_index <= 5445)) || ((pixel_index >= 5450) && (pixel_index <= 5451)) || ((pixel_index >= 5460) && (pixel_index <= 5461)) || ((pixel_index >= 5504) && (pixel_index <= 5506)) || ((pixel_index >= 5514) && (pixel_index <= 5515)) || ((pixel_index >= 5524) && (pixel_index <= 5525)) || ((pixel_index >= 5536) && (pixel_index <= 5537)) || ((pixel_index >= 5540) && (pixel_index <= 5541)) || ((pixel_index >= 5546) && (pixel_index <= 5547)) || ((pixel_index >= 5556) && (pixel_index <= 5557)) || ((pixel_index >= 5599) && (pixel_index <= 5601)) || ((pixel_index >= 5610) && (pixel_index <= 5617)) || ((pixel_index >= 5620) && (pixel_index <= 5627)) || ((pixel_index >= 5634) && (pixel_index <= 5635)) || ((pixel_index >= 5642) && (pixel_index <= 5649)) || ((pixel_index >= 5652) && (pixel_index <= 5659)) || ((pixel_index >= 5695) && (pixel_index <= 5696)) || ((pixel_index >= 5706) && (pixel_index <= 5713)) || ((pixel_index >= 5716) && (pixel_index <= 5723)) || ((pixel_index >= 5730) && (pixel_index <= 5731)) || ((pixel_index >= 5738) && (pixel_index <= 5745)) || (pixel_index >= 5748) && (pixel_index <= 5755)) oled_data = 16'b1111111111111111;
            else if (((pixel_index >= 628) && (pixel_index <= 629)) || ((pixel_index >= 636) && (pixel_index <= 637)) || ((pixel_index >= 640) && (pixel_index <= 645)) || ((pixel_index >= 648) && (pixel_index <= 649)) || ((pixel_index >= 654) && (pixel_index <= 655)) || ((pixel_index >= 724) && (pixel_index <= 725)) || pixel_index == 733 || ((pixel_index >= 736) && (pixel_index <= 737)) || ((pixel_index >= 739) && (pixel_index <= 740)) || ((pixel_index >= 744) && (pixel_index <= 745)) || ((pixel_index >= 750) && (pixel_index <= 751)) || ((pixel_index >= 820) && (pixel_index <= 821)) || ((pixel_index >= 828) && (pixel_index <= 829)) || ((pixel_index >= 834) && (pixel_index <= 835)) || ((pixel_index >= 840) && (pixel_index <= 843)) || ((pixel_index >= 846) && (pixel_index <= 847)) || pixel_index == 917 || ((pixel_index >= 924) && (pixel_index <= 925)) || ((pixel_index >= 930) && (pixel_index <= 931)) || ((pixel_index >= 936) && (pixel_index <= 937)) || pixel_index == 939 || ((pixel_index >= 942) && (pixel_index <= 943)) || ((pixel_index >= 1012) && (pixel_index <= 1013)) || ((pixel_index >= 1016) && (pixel_index <= 1017)) || ((pixel_index >= 1020) && (pixel_index <= 1021)) || ((pixel_index >= 1026) && (pixel_index <= 1027)) || ((pixel_index >= 1032) && (pixel_index <= 1033)) || ((pixel_index >= 1036) && (pixel_index <= 1037)) || pixel_index == 1039 || ((pixel_index >= 1108) && (pixel_index <= 1109)) || ((pixel_index >= 1112) && (pixel_index <= 1113)) || ((pixel_index >= 1116) && (pixel_index <= 1117)) || pixel_index == 1123 || pixel_index == 1128 || ((pixel_index >= 1132) && (pixel_index <= 1135)) || pixel_index == 1204 || ((pixel_index >= 1206) && (pixel_index <= 1207)) || ((pixel_index >= 1210) && (pixel_index <= 1211)) || pixel_index == 1213 || ((pixel_index >= 1218) && (pixel_index <= 1219)) || ((pixel_index >= 1224) && (pixel_index <= 1225)) || ((pixel_index >= 1230) && (pixel_index <= 1231)) || ((pixel_index >= 1300) && (pixel_index <= 1303)) || ((pixel_index >= 1307) && (pixel_index <= 1309)) || ((pixel_index >= 1314) && (pixel_index <= 1315)) || ((pixel_index >= 1320) && (pixel_index <= 1321)) || ((pixel_index >= 1326) && (pixel_index <= 1327)) || ((pixel_index >= 1396) && (pixel_index <= 1397)) || ((pixel_index >= 1404) && (pixel_index <= 1405)) || ((pixel_index >= 1408) && (pixel_index <= 1413)) || pixel_index == 1416 || ((pixel_index >= 1422) && (pixel_index <= 1423)) || ((pixel_index >= 1492) && (pixel_index <= 1493)) || ((pixel_index >= 1500) && (pixel_index <= 1501)) || pixel_index == 1504 || pixel_index == 1506 || ((pixel_index >= 1508) && (pixel_index <= 1509)) || ((pixel_index >= 1512) && (pixel_index <= 1513)) || (pixel_index >= 1518) && (pixel_index <= 1519) || pixel_index == 732 || pixel_index == 738 || pixel_index == 741 || pixel_index == 916 || pixel_index == 938 || pixel_index == 1038 || pixel_index == 1122 || pixel_index == 1129 || pixel_index == 1205 || pixel_index == 1212 || pixel_index == 1306 || pixel_index == 1417 || pixel_index == 1505 || pixel_index == 1507) oled_data = 16'b0001011101111111;
            else oled_data = 16'b0000000001000100;
        end
        else if (result == 2'b10) begin // player lose
            if (((pixel_index >= 194) && (pixel_index <= 285)) || ((pixel_index >= 290) && (pixel_index <= 381)) || ((pixel_index >= 386) && (pixel_index <= 387)) || ((pixel_index >= 476) && (pixel_index <= 477)) || ((pixel_index >= 482) && (pixel_index <= 483)) || ((pixel_index >= 572) && (pixel_index <= 573)) || ((pixel_index >= 578) && (pixel_index <= 579)) || ((pixel_index >= 587) && (pixel_index <= 588)) || ((pixel_index >= 595) && (pixel_index <= 596)) || ((pixel_index >= 601) && (pixel_index <= 604)) || ((pixel_index >= 609) && (pixel_index <= 610)) || ((pixel_index >= 615) && (pixel_index <= 616)) || ((pixel_index >= 668) && (pixel_index <= 669)) || ((pixel_index >= 674) && (pixel_index <= 675)) || ((pixel_index >= 683) && (pixel_index <= 684)) || ((pixel_index >= 691) && (pixel_index <= 692)) || ((pixel_index >= 697) && (pixel_index <= 700)) || ((pixel_index >= 705) && (pixel_index <= 706)) || ((pixel_index >= 711) && (pixel_index <= 712)) || ((pixel_index >= 764) && (pixel_index <= 765)) || ((pixel_index >= 770) && (pixel_index <= 771)) || ((pixel_index >= 779) && (pixel_index <= 780)) || ((pixel_index >= 787) && (pixel_index <= 788)) || ((pixel_index >= 791) && (pixel_index <= 792)) || ((pixel_index >= 797) && (pixel_index <= 798)) || ((pixel_index >= 801) && (pixel_index <= 802)) || ((pixel_index >= 807) && (pixel_index <= 808)) || ((pixel_index >= 860) && (pixel_index <= 861)) || ((pixel_index >= 866) && (pixel_index <= 867)) || ((pixel_index >= 875) && (pixel_index <= 876)) || ((pixel_index >= 883) && (pixel_index <= 884)) || ((pixel_index >= 887) && (pixel_index <= 888)) || ((pixel_index >= 893) && (pixel_index <= 894)) || ((pixel_index >= 897) && (pixel_index <= 898)) || ((pixel_index >= 903) && (pixel_index <= 904)) || ((pixel_index >= 956) && (pixel_index <= 957)) || ((pixel_index >= 962) && (pixel_index <= 963)) || ((pixel_index >= 973) && (pixel_index <= 978)) || ((pixel_index >= 983) && (pixel_index <= 984)) || ((pixel_index >= 989) && (pixel_index <= 990)) || ((pixel_index >= 993) && (pixel_index <= 994)) || ((pixel_index >= 999) && (pixel_index <= 1000)) || ((pixel_index >= 1052) && (pixel_index <= 1053)) || ((pixel_index >= 1058) && (pixel_index <= 1059)) || ((pixel_index >= 1069) && (pixel_index <= 1074)) || ((pixel_index >= 1079) && (pixel_index <= 1080)) || ((pixel_index >= 1085) && (pixel_index <= 1086)) || ((pixel_index >= 1089) && (pixel_index <= 1090)) || ((pixel_index >= 1095) && (pixel_index <= 1096)) || ((pixel_index >= 1148) && (pixel_index <= 1149)) || ((pixel_index >= 1154) && (pixel_index <= 1155)) || ((pixel_index >= 1167) && (pixel_index <= 1168)) || ((pixel_index >= 1175) && (pixel_index <= 1176)) || ((pixel_index >= 1181) && (pixel_index <= 1182)) || ((pixel_index >= 1185) && (pixel_index <= 1186)) || ((pixel_index >= 1191) && (pixel_index <= 1192)) || ((pixel_index >= 1244) && (pixel_index <= 1245)) || ((pixel_index >= 1250) && (pixel_index <= 1251)) || ((pixel_index >= 1263) && (pixel_index <= 1264)) || ((pixel_index >= 1271) && (pixel_index <= 1272)) || ((pixel_index >= 1277) && (pixel_index <= 1278)) || ((pixel_index >= 1281) && (pixel_index <= 1282)) || ((pixel_index >= 1287) && (pixel_index <= 1288)) || ((pixel_index >= 1340) && (pixel_index <= 1341)) || ((pixel_index >= 1346) && (pixel_index <= 1347)) || ((pixel_index >= 1359) && (pixel_index <= 1360)) || ((pixel_index >= 1369) && (pixel_index <= 1372)) || ((pixel_index >= 1379) && (pixel_index <= 1382)) || ((pixel_index >= 1436) && (pixel_index <= 1437)) || ((pixel_index >= 1442) && (pixel_index <= 1443)) || ((pixel_index >= 1455) && (pixel_index <= 1456)) || ((pixel_index >= 1465) && (pixel_index <= 1468)) || ((pixel_index >= 1475) && (pixel_index <= 1478)) || ((pixel_index >= 1532) && (pixel_index <= 1533)) || ((pixel_index >= 1538) && (pixel_index <= 1539)) || ((pixel_index >= 1628) && (pixel_index <= 1629)) || ((pixel_index >= 1634) && (pixel_index <= 1635)) || ((pixel_index >= 1724) && (pixel_index <= 1725)) || ((pixel_index >= 1730) && (pixel_index <= 1821)) || ((pixel_index >= 1826) && (pixel_index <= 1917)) || ((pixel_index >= 3676) && (pixel_index <= 3681)) || ((pixel_index >= 3688) && (pixel_index <= 3691)) || ((pixel_index >= 3698) && (pixel_index <= 3701)) || ((pixel_index >= 3706) && (pixel_index <= 3707)) || ((pixel_index >= 3712) && (pixel_index <= 3713)) || ((pixel_index >= 3720) && (pixel_index <= 3729)) || ((pixel_index >= 3734) && (pixel_index <= 3737)) || ((pixel_index >= 3772) && (pixel_index <= 3777)) || ((pixel_index >= 3784) && (pixel_index <= 3787)) || ((pixel_index >= 3794) && (pixel_index <= 3797)) || ((pixel_index >= 3802) && (pixel_index <= 3803)) || ((pixel_index >= 3808) && (pixel_index <= 3809)) || ((pixel_index >= 3816) && (pixel_index <= 3825)) || ((pixel_index >= 3830) && (pixel_index <= 3833)) || ((pixel_index >= 3868) && (pixel_index <= 3869)) || ((pixel_index >= 3874) && (pixel_index <= 3875)) || ((pixel_index >= 3878) && (pixel_index <= 3879)) || ((pixel_index >= 3884) && (pixel_index <= 3885)) || ((pixel_index >= 3888) && (pixel_index <= 3889)) || ((pixel_index >= 3894) && (pixel_index <= 3895)) || ((pixel_index >= 3898) && (pixel_index <= 3899)) || ((pixel_index >= 3902) && (pixel_index <= 3903)) || ((pixel_index >= 3916) && (pixel_index <= 3917)) || ((pixel_index >= 3924) && (pixel_index <= 3925)) || ((pixel_index >= 3930) && (pixel_index <= 3931)) || ((pixel_index >= 3964) && (pixel_index <= 3965)) || ((pixel_index >= 3970) && (pixel_index <= 3971)) || ((pixel_index >= 3974) && (pixel_index <= 3975)) || ((pixel_index >= 3980) && (pixel_index <= 3981)) || ((pixel_index >= 3984) && (pixel_index <= 3985)) || ((pixel_index >= 3990) && (pixel_index <= 3991)) || ((pixel_index >= 3994) && (pixel_index <= 3995)) || ((pixel_index >= 3998) && (pixel_index <= 3999)) || ((pixel_index >= 4012) && (pixel_index <= 4013)) || ((pixel_index >= 4020) && (pixel_index <= 4021)) || ((pixel_index >= 4026) && (pixel_index <= 4027)) || ((pixel_index >= 4060) && (pixel_index <= 4065)) || ((pixel_index >= 4070) && (pixel_index <= 4077)) || ((pixel_index >= 4080) && (pixel_index <= 4081)) || ((pixel_index >= 4090) && (pixel_index <= 4093)) || ((pixel_index >= 4108) && (pixel_index <= 4109)) || ((pixel_index >= 4116) && (pixel_index <= 4117)) || ((pixel_index >= 4122) && (pixel_index <= 4123)) || ((pixel_index >= 4156) && (pixel_index <= 4161)) || ((pixel_index >= 4166) && (pixel_index <= 4173)) || ((pixel_index >= 4176) && (pixel_index <= 4177)) || ((pixel_index >= 4186) && (pixel_index <= 4189)) || ((pixel_index >= 4204) && (pixel_index <= 4205)) || ((pixel_index >= 4212) && (pixel_index <= 4213)) || ((pixel_index >= 4218) && (pixel_index <= 4219)) || ((pixel_index >= 4252) && (pixel_index <= 4253)) || ((pixel_index >= 4258) && (pixel_index <= 4259)) || ((pixel_index >= 4262) && (pixel_index <= 4263)) || ((pixel_index >= 4268) && (pixel_index <= 4269)) || ((pixel_index >= 4272) && (pixel_index <= 4273)) || ((pixel_index >= 4278) && (pixel_index <= 4279)) || ((pixel_index >= 4282) && (pixel_index <= 4283)) || ((pixel_index >= 4286) && (pixel_index <= 4287)) || ((pixel_index >= 4300) && (pixel_index <= 4301)) || ((pixel_index >= 4308) && (pixel_index <= 4309)) || ((pixel_index >= 4314) && (pixel_index <= 4315)) || ((pixel_index >= 4348) && (pixel_index <= 4349)) || ((pixel_index >= 4354) && (pixel_index <= 4355)) || ((pixel_index >= 4358) && (pixel_index <= 4359)) || ((pixel_index >= 4364) && (pixel_index <= 4365)) || ((pixel_index >= 4368) && (pixel_index <= 4369)) || ((pixel_index >= 4374) && (pixel_index <= 4375)) || ((pixel_index >= 4378) && (pixel_index <= 4379)) || ((pixel_index >= 4382) && (pixel_index <= 4383)) || ((pixel_index >= 4396) && (pixel_index <= 4397)) || ((pixel_index >= 4404) && (pixel_index <= 4405)) || ((pixel_index >= 4410) && (pixel_index <= 4411)) || ((pixel_index >= 4444) && (pixel_index <= 4449)) || ((pixel_index >= 4454) && (pixel_index <= 4455)) || ((pixel_index >= 4460) && (pixel_index <= 4461)) || ((pixel_index >= 4466) && (pixel_index <= 4469)) || ((pixel_index >= 4474) && (pixel_index <= 4475)) || ((pixel_index >= 4480) && (pixel_index <= 4481)) || ((pixel_index >= 4492) && (pixel_index <= 4493)) || ((pixel_index >= 4502) && (pixel_index <= 4505)) || ((pixel_index >= 4540) && (pixel_index <= 4545)) || ((pixel_index >= 4550) && (pixel_index <= 4551)) || ((pixel_index >= 4556) && (pixel_index <= 4557)) || ((pixel_index >= 4562) && (pixel_index <= 4565)) || ((pixel_index >= 4570) && (pixel_index <= 4571)) || ((pixel_index >= 4576) && (pixel_index <= 4577)) || ((pixel_index >= 4588) && (pixel_index <= 4589)) || ((pixel_index >= 4598) && (pixel_index <= 4601)) || ((pixel_index >= 4819) && (pixel_index <= 4820)) || ((pixel_index >= 4830) && (pixel_index <= 4831)) || ((pixel_index >= 4840) && (pixel_index <= 4847)) || ((pixel_index >= 4850) && (pixel_index <= 4851)) || ((pixel_index >= 4858) && (pixel_index <= 4859)) || ((pixel_index >= 4862) && (pixel_index <= 4869)) || ((pixel_index >= 4872) && (pixel_index <= 4873)) || ((pixel_index >= 4888) && (pixel_index <= 4889)) || ((pixel_index >= 4915) && (pixel_index <= 4917)) || ((pixel_index >= 4926) && (pixel_index <= 4927)) || ((pixel_index >= 4936) && (pixel_index <= 4943)) || ((pixel_index >= 4946) && (pixel_index <= 4947)) || ((pixel_index >= 4954) && (pixel_index <= 4955)) || ((pixel_index >= 4958) && (pixel_index <= 4965)) || ((pixel_index >= 4968) && (pixel_index <= 4969)) || ((pixel_index >= 4984) && (pixel_index <= 4985)) || ((pixel_index >= 5012) && (pixel_index <= 5014)) || ((pixel_index >= 5022) && (pixel_index <= 5023)) || ((pixel_index >= 5032) && (pixel_index <= 5033)) || ((pixel_index >= 5042) && (pixel_index <= 5043)) || ((pixel_index >= 5050) && (pixel_index <= 5051)) || ((pixel_index >= 5054) && (pixel_index <= 5055)) || ((pixel_index >= 5064) && (pixel_index <= 5065)) || ((pixel_index >= 5078) && (pixel_index <= 5081)) || ((pixel_index >= 5109) && (pixel_index <= 5111)) || ((pixel_index >= 5118) && (pixel_index <= 5119)) || ((pixel_index >= 5128) && (pixel_index <= 5129)) || ((pixel_index >= 5138) && (pixel_index <= 5139)) || ((pixel_index >= 5146) && (pixel_index <= 5147)) || ((pixel_index >= 5150) && (pixel_index <= 5151)) || ((pixel_index >= 5160) && (pixel_index <= 5161)) || ((pixel_index >= 5174) && (pixel_index <= 5177)) || ((pixel_index >= 5193) && (pixel_index <= 5208)) || ((pixel_index >= 5214) && (pixel_index <= 5215)) || ((pixel_index >= 5224) && (pixel_index <= 5229)) || ((pixel_index >= 5236) && (pixel_index <= 5237)) || ((pixel_index >= 5240) && (pixel_index <= 5241)) || ((pixel_index >= 5246) && (pixel_index <= 5251)) || ((pixel_index >= 5256) && (pixel_index <= 5257)) || ((pixel_index >= 5272) && (pixel_index <= 5273)) || ((pixel_index >= 5289) && (pixel_index <= 5304)) || ((pixel_index >= 5310) && (pixel_index <= 5311)) || ((pixel_index >= 5320) && (pixel_index <= 5325)) || ((pixel_index >= 5332) && (pixel_index <= 5333)) || ((pixel_index >= 5336) && (pixel_index <= 5337)) || ((pixel_index >= 5342) && (pixel_index <= 5347)) || ((pixel_index >= 5352) && (pixel_index <= 5353)) || ((pixel_index >= 5368) && (pixel_index <= 5369)) || ((pixel_index >= 5397) && (pixel_index <= 5399)) || ((pixel_index >= 5406) && (pixel_index <= 5407)) || ((pixel_index >= 5416) && (pixel_index <= 5417)) || ((pixel_index >= 5428) && (pixel_index <= 5429)) || ((pixel_index >= 5432) && (pixel_index <= 5433)) || ((pixel_index >= 5438) && (pixel_index <= 5439)) || ((pixel_index >= 5448) && (pixel_index <= 5449)) || ((pixel_index >= 5464) && (pixel_index <= 5465)) || ((pixel_index >= 5492) && (pixel_index <= 5494)) || ((pixel_index >= 5502) && (pixel_index <= 5503)) || ((pixel_index >= 5512) && (pixel_index <= 5513)) || ((pixel_index >= 5524) && (pixel_index <= 5525)) || ((pixel_index >= 5528) && (pixel_index <= 5529)) || ((pixel_index >= 5534) && (pixel_index <= 5535)) || ((pixel_index >= 5544) && (pixel_index <= 5545)) || ((pixel_index >= 5560) && (pixel_index <= 5561)) || ((pixel_index >= 5587) && (pixel_index <= 5589)) || ((pixel_index >= 5598) && (pixel_index <= 5605)) || ((pixel_index >= 5608) && (pixel_index <= 5615)) || ((pixel_index >= 5622) && (pixel_index <= 5623)) || ((pixel_index >= 5630) && (pixel_index <= 5637)) || ((pixel_index >= 5640) && (pixel_index <= 5647)) || ((pixel_index >= 5654) && (pixel_index <= 5659)) || ((pixel_index >= 5683) && (pixel_index <= 5684)) || ((pixel_index >= 5694) && (pixel_index <= 5701)) || ((pixel_index >= 5704) && (pixel_index <= 5711)) || ((pixel_index >= 5718) && (pixel_index <= 5719)) || ((pixel_index >= 5726) && (pixel_index <= 5733)) || ((pixel_index >= 5736) && (pixel_index <= 5743)) || (pixel_index >= 5750) && (pixel_index <= 5755)) oled_data = 16'b1111111111111111;
            else if (((pixel_index >= 623) && (pixel_index <= 624)) || pixel_index == 635 || ((pixel_index >= 637) && (pixel_index <= 638)) || ((pixel_index >= 645) && (pixel_index <= 650)) || ((pixel_index >= 653) && (pixel_index <= 659)) || ((pixel_index >= 719) && (pixel_index <= 720)) || ((pixel_index >= 731) && (pixel_index <= 732)) || pixel_index == 734 || pixel_index == 741 || pixel_index == 743 || pixel_index == 745 || pixel_index == 749 || pixel_index == 751 || pixel_index == 753 || ((pixel_index >= 755) && (pixel_index <= 756)) || pixel_index == 815 || ((pixel_index >= 825) && (pixel_index <= 826)) || ((pixel_index >= 831) && (pixel_index <= 832)) || pixel_index == 835 || pixel_index == 845 || ((pixel_index >= 911) && (pixel_index <= 912)) || pixel_index == 921 || pixel_index == 928 || ((pixel_index >= 931) && (pixel_index <= 932)) || pixel_index == 942 || pixel_index == 1007 || ((pixel_index >= 1017) && (pixel_index <= 1018)) || pixel_index == 1023 || ((pixel_index >= 1029) && (pixel_index <= 1032)) || pixel_index == 1037 || ((pixel_index >= 1039) && (pixel_index <= 1042)) || ((pixel_index >= 1103) && (pixel_index <= 1104)) || pixel_index == 1114 || ((pixel_index >= 1119) && (pixel_index <= 1120)) || pixel_index == 1126 || pixel_index == 1128 || pixel_index == 1133 || pixel_index == 1135 || pixel_index == 1138 || pixel_index == 1199 || pixel_index == 1209 || pixel_index == 1215 || ((pixel_index >= 1225) && (pixel_index <= 1226)) || ((pixel_index >= 1229) && (pixel_index <= 1230)) || ((pixel_index >= 1295) && (pixel_index <= 1296)) || ((pixel_index >= 1305) && (pixel_index <= 1306)) || ((pixel_index >= 1311) && (pixel_index <= 1312)) || pixel_index == 1322 || pixel_index == 1326 || pixel_index == 1391 || ((pixel_index >= 1393) && (pixel_index <= 1396)) || pixel_index == 1398 || ((pixel_index >= 1403) && (pixel_index <= 1406)) || ((pixel_index >= 1411) && (pixel_index <= 1416)) || pixel_index == 1421 || ((pixel_index >= 1423) && (pixel_index <= 1428)) || ((pixel_index >= 1487) && (pixel_index <= 1488)) || pixel_index == 1490 || ((pixel_index >= 1492) && (pixel_index <= 1493)) || pixel_index == 1500 || pixel_index == 1507 || pixel_index == 1512 || ((pixel_index >= 1517) && (pixel_index <= 1518)) || pixel_index == 1521 || pixel_index == 1524 || pixel_index == 636 || pixel_index == 660 || pixel_index == 733 || pixel_index == 742 || pixel_index == 746 || pixel_index == 750 || pixel_index == 752 || pixel_index == 754 || pixel_index == 816 || pixel_index == 836 || pixel_index == 846 || pixel_index == 922 || pixel_index == 927 || pixel_index == 1008 || pixel_index == 1024 || pixel_index == 1038 || pixel_index == 1113 || pixel_index == 1125 || pixel_index == 1127 || pixel_index == 1134 || ((pixel_index >= 1136) && (pixel_index <= 1137)) || pixel_index == 1200 || pixel_index == 1210 || pixel_index == 1216 || pixel_index == 1321 || pixel_index == 1392 || pixel_index == 1397 || pixel_index == 1422 || pixel_index == 1489 || pixel_index == 1491 || pixel_index == 1494 || pixel_index == 1499 || ((pixel_index >= 1501) && (pixel_index <= 1502)) || pixel_index == 1508 || ((pixel_index >= 1510) && (pixel_index <= 1511)) || ((pixel_index >= 1519) && (pixel_index <= 1520)) || pixel_index == 1522 || pixel_index == 744 || pixel_index == 1325 || pixel_index == 1523 || pixel_index == 941 || pixel_index == 1509) oled_data = 16'b1111100001011000;
            else oled_data = 16'b0000000001000100;
        end
        else if (result == 2'b11) begin // draw
            if (((pixel_index >= 194) && (pixel_index <= 285)) || ((pixel_index >= 290) && (pixel_index <= 381)) || ((pixel_index >= 386) && (pixel_index <= 387)) || ((pixel_index >= 476) && (pixel_index <= 477)) || ((pixel_index >= 482) && (pixel_index <= 483)) || ((pixel_index >= 572) && (pixel_index <= 573)) || ((pixel_index >= 578) && (pixel_index <= 579)) || ((pixel_index >= 604) && (pixel_index <= 609)) || ((pixel_index >= 614) && (pixel_index <= 619)) || ((pixel_index >= 626) && (pixel_index <= 629)) || ((pixel_index >= 634) && (pixel_index <= 635)) || ((pixel_index >= 642) && (pixel_index <= 643)) || ((pixel_index >= 668) && (pixel_index <= 669)) || ((pixel_index >= 674) && (pixel_index <= 675)) || ((pixel_index >= 700) && (pixel_index <= 705)) || ((pixel_index >= 710) && (pixel_index <= 715)) || ((pixel_index >= 722) && (pixel_index <= 725)) || ((pixel_index >= 730) && (pixel_index <= 731)) || ((pixel_index >= 738) && (pixel_index <= 739)) || ((pixel_index >= 764) && (pixel_index <= 765)) || ((pixel_index >= 770) && (pixel_index <= 771)) || ((pixel_index >= 796) && (pixel_index <= 797)) || ((pixel_index >= 802) && (pixel_index <= 803)) || ((pixel_index >= 806) && (pixel_index <= 807)) || ((pixel_index >= 812) && (pixel_index <= 813)) || ((pixel_index >= 816) && (pixel_index <= 817)) || ((pixel_index >= 822) && (pixel_index <= 823)) || ((pixel_index >= 826) && (pixel_index <= 827)) || ((pixel_index >= 834) && (pixel_index <= 835)) || ((pixel_index >= 860) && (pixel_index <= 861)) || ((pixel_index >= 866) && (pixel_index <= 867)) || ((pixel_index >= 892) && (pixel_index <= 893)) || ((pixel_index >= 898) && (pixel_index <= 899)) || ((pixel_index >= 902) && (pixel_index <= 903)) || ((pixel_index >= 908) && (pixel_index <= 909)) || ((pixel_index >= 912) && (pixel_index <= 913)) || ((pixel_index >= 918) && (pixel_index <= 919)) || ((pixel_index >= 922) && (pixel_index <= 923)) || ((pixel_index >= 930) && (pixel_index <= 931)) || ((pixel_index >= 956) && (pixel_index <= 957)) || ((pixel_index >= 962) && (pixel_index <= 963)) || ((pixel_index >= 988) && (pixel_index <= 989)) || ((pixel_index >= 994) && (pixel_index <= 995)) || ((pixel_index >= 998) && (pixel_index <= 1003)) || ((pixel_index >= 1008) && (pixel_index <= 1015)) || ((pixel_index >= 1018) && (pixel_index <= 1019)) || ((pixel_index >= 1022) && (pixel_index <= 1023)) || ((pixel_index >= 1026) && (pixel_index <= 1027)) || ((pixel_index >= 1052) && (pixel_index <= 1053)) || ((pixel_index >= 1058) && (pixel_index <= 1059)) || ((pixel_index >= 1084) && (pixel_index <= 1085)) || ((pixel_index >= 1090) && (pixel_index <= 1091)) || ((pixel_index >= 1094) && (pixel_index <= 1099)) || ((pixel_index >= 1104) && (pixel_index <= 1111)) || ((pixel_index >= 1114) && (pixel_index <= 1115)) || ((pixel_index >= 1118) && (pixel_index <= 1119)) || ((pixel_index >= 1122) && (pixel_index <= 1123)) || ((pixel_index >= 1148) && (pixel_index <= 1149)) || ((pixel_index >= 1154) && (pixel_index <= 1155)) || ((pixel_index >= 1180) && (pixel_index <= 1181)) || ((pixel_index >= 1186) && (pixel_index <= 1187)) || ((pixel_index >= 1190) && (pixel_index <= 1191)) || ((pixel_index >= 1194) && (pixel_index <= 1195)) || ((pixel_index >= 1200) && (pixel_index <= 1201)) || ((pixel_index >= 1206) && (pixel_index <= 1207)) || ((pixel_index >= 1210) && (pixel_index <= 1213)) || ((pixel_index >= 1216) && (pixel_index <= 1219)) || ((pixel_index >= 1244) && (pixel_index <= 1245)) || ((pixel_index >= 1250) && (pixel_index <= 1251)) || ((pixel_index >= 1276) && (pixel_index <= 1277)) || ((pixel_index >= 1282) && (pixel_index <= 1283)) || ((pixel_index >= 1286) && (pixel_index <= 1287)) || ((pixel_index >= 1290) && (pixel_index <= 1291)) || ((pixel_index >= 1296) && (pixel_index <= 1297)) || ((pixel_index >= 1302) && (pixel_index <= 1303)) || ((pixel_index >= 1306) && (pixel_index <= 1309)) || ((pixel_index >= 1312) && (pixel_index <= 1315)) || ((pixel_index >= 1340) && (pixel_index <= 1341)) || ((pixel_index >= 1346) && (pixel_index <= 1347)) || ((pixel_index >= 1372) && (pixel_index <= 1377)) || ((pixel_index >= 1382) && (pixel_index <= 1383)) || ((pixel_index >= 1388) && (pixel_index <= 1389)) || ((pixel_index >= 1392) && (pixel_index <= 1393)) || ((pixel_index >= 1398) && (pixel_index <= 1399)) || ((pixel_index >= 1402) && (pixel_index <= 1403)) || ((pixel_index >= 1410) && (pixel_index <= 1411)) || ((pixel_index >= 1436) && (pixel_index <= 1437)) || ((pixel_index >= 1442) && (pixel_index <= 1443)) || ((pixel_index >= 1468) && (pixel_index <= 1473)) || ((pixel_index >= 1478) && (pixel_index <= 1479)) || ((pixel_index >= 1484) && (pixel_index <= 1485)) || ((pixel_index >= 1488) && (pixel_index <= 1489)) || ((pixel_index >= 1494) && (pixel_index <= 1495)) || ((pixel_index >= 1498) && (pixel_index <= 1499)) || ((pixel_index >= 1506) && (pixel_index <= 1507)) || ((pixel_index >= 1532) && (pixel_index <= 1533)) || ((pixel_index >= 1538) && (pixel_index <= 1539)) || ((pixel_index >= 1628) && (pixel_index <= 1629)) || ((pixel_index >= 1634) && (pixel_index <= 1635)) || ((pixel_index >= 1724) && (pixel_index <= 1725)) || ((pixel_index >= 1730) && (pixel_index <= 1821)) || ((pixel_index >= 1826) && (pixel_index <= 1917)) || ((pixel_index >= 3668) && (pixel_index <= 3673)) || ((pixel_index >= 3678) && (pixel_index <= 3685)) || ((pixel_index >= 3690) && (pixel_index <= 3695)) || ((pixel_index >= 3698) && (pixel_index <= 3707)) || ((pixel_index >= 3712) && (pixel_index <= 3715)) || ((pixel_index >= 3720) && (pixel_index <= 3725)) || ((pixel_index >= 3730) && (pixel_index <= 3739)) || ((pixel_index >= 3764) && (pixel_index <= 3769)) || ((pixel_index >= 3774) && (pixel_index <= 3781)) || ((pixel_index >= 3786) && (pixel_index <= 3791)) || ((pixel_index >= 3794) && (pixel_index <= 3803)) || ((pixel_index >= 3808) && (pixel_index <= 3811)) || ((pixel_index >= 3816) && (pixel_index <= 3821)) || ((pixel_index >= 3826) && (pixel_index <= 3835)) || ((pixel_index >= 3860) && (pixel_index <= 3861)) || ((pixel_index >= 3866) && (pixel_index <= 3867)) || ((pixel_index >= 3870) && (pixel_index <= 3871)) || ((pixel_index >= 3880) && (pixel_index <= 3881)) || ((pixel_index >= 3894) && (pixel_index <= 3895)) || ((pixel_index >= 3902) && (pixel_index <= 3903)) || ((pixel_index >= 3908) && (pixel_index <= 3909)) || ((pixel_index >= 3912) && (pixel_index <= 3913)) || ((pixel_index >= 3918) && (pixel_index <= 3919)) || ((pixel_index >= 3926) && (pixel_index <= 3927)) || ((pixel_index >= 3956) && (pixel_index <= 3957)) || ((pixel_index >= 3962) && (pixel_index <= 3963)) || ((pixel_index >= 3966) && (pixel_index <= 3967)) || ((pixel_index >= 3976) && (pixel_index <= 3977)) || ((pixel_index >= 3990) && (pixel_index <= 3991)) || ((pixel_index >= 3998) && (pixel_index <= 3999)) || ((pixel_index >= 4004) && (pixel_index <= 4005)) || ((pixel_index >= 4008) && (pixel_index <= 4009)) || ((pixel_index >= 4014) && (pixel_index <= 4015)) || ((pixel_index >= 4022) && (pixel_index <= 4023)) || ((pixel_index >= 4052) && (pixel_index <= 4057)) || ((pixel_index >= 4062) && (pixel_index <= 4067)) || ((pixel_index >= 4074) && (pixel_index <= 4077)) || ((pixel_index >= 4086) && (pixel_index <= 4087)) || ((pixel_index >= 4094) && (pixel_index <= 4101)) || ((pixel_index >= 4104) && (pixel_index <= 4109)) || ((pixel_index >= 4118) && (pixel_index <= 4119)) || ((pixel_index >= 4148) && (pixel_index <= 4153)) || ((pixel_index >= 4158) && (pixel_index <= 4163)) || ((pixel_index >= 4170) && (pixel_index <= 4173)) || ((pixel_index >= 4182) && (pixel_index <= 4183)) || ((pixel_index >= 4190) && (pixel_index <= 4197)) || ((pixel_index >= 4200) && (pixel_index <= 4205)) || ((pixel_index >= 4214) && (pixel_index <= 4215)) || ((pixel_index >= 4244) && (pixel_index <= 4245)) || ((pixel_index >= 4248) && (pixel_index <= 4249)) || ((pixel_index >= 4254) && (pixel_index <= 4255)) || ((pixel_index >= 4270) && (pixel_index <= 4271)) || ((pixel_index >= 4278) && (pixel_index <= 4279)) || ((pixel_index >= 4286) && (pixel_index <= 4287)) || ((pixel_index >= 4292) && (pixel_index <= 4293)) || ((pixel_index >= 4296) && (pixel_index <= 4297)) || ((pixel_index >= 4300) && (pixel_index <= 4301)) || ((pixel_index >= 4310) && (pixel_index <= 4311)) || ((pixel_index >= 4340) && (pixel_index <= 4341)) || ((pixel_index >= 4344) && (pixel_index <= 4345)) || ((pixel_index >= 4350) && (pixel_index <= 4351)) || ((pixel_index >= 4366) && (pixel_index <= 4367)) || ((pixel_index >= 4374) && (pixel_index <= 4375)) || ((pixel_index >= 4382) && (pixel_index <= 4383)) || ((pixel_index >= 4388) && (pixel_index <= 4389)) || ((pixel_index >= 4392) && (pixel_index <= 4393)) || ((pixel_index >= 4396) && (pixel_index <= 4397)) || ((pixel_index >= 4406) && (pixel_index <= 4407)) || ((pixel_index >= 4436) && (pixel_index <= 4437)) || ((pixel_index >= 4442) && (pixel_index <= 4443)) || ((pixel_index >= 4446) && (pixel_index <= 4453)) || ((pixel_index >= 4456) && (pixel_index <= 4461)) || ((pixel_index >= 4470) && (pixel_index <= 4471)) || ((pixel_index >= 4478) && (pixel_index <= 4479)) || ((pixel_index >= 4484) && (pixel_index <= 4485)) || ((pixel_index >= 4488) && (pixel_index <= 4489)) || ((pixel_index >= 4494) && (pixel_index <= 4495)) || ((pixel_index >= 4502) && (pixel_index <= 4503)) || ((pixel_index >= 4532) && (pixel_index <= 4533)) || ((pixel_index >= 4538) && (pixel_index <= 4539)) || ((pixel_index >= 4542) && (pixel_index <= 4549)) || ((pixel_index >= 4552) && (pixel_index <= 4557)) || ((pixel_index >= 4566) && (pixel_index <= 4567)) || ((pixel_index >= 4574) && (pixel_index <= 4575)) || ((pixel_index >= 4580) && (pixel_index <= 4581)) || ((pixel_index >= 4584) && (pixel_index <= 4585)) || ((pixel_index >= 4590) && (pixel_index <= 4591)) || ((pixel_index >= 4598) && (pixel_index <= 4599)) || ((pixel_index >= 4831) && (pixel_index <= 4832)) || ((pixel_index >= 4842) && (pixel_index <= 4843)) || ((pixel_index >= 4852) && (pixel_index <= 4859)) || ((pixel_index >= 4862) && (pixel_index <= 4863)) || ((pixel_index >= 4870) && (pixel_index <= 4871)) || ((pixel_index >= 4874) && (pixel_index <= 4881)) || ((pixel_index >= 4884) && (pixel_index <= 4885)) || ((pixel_index >= 4927) && (pixel_index <= 4929)) || ((pixel_index >= 4938) && (pixel_index <= 4939)) || ((pixel_index >= 4948) && (pixel_index <= 4955)) || ((pixel_index >= 4958) && (pixel_index <= 4959)) || ((pixel_index >= 4966) && (pixel_index <= 4967)) || ((pixel_index >= 4970) && (pixel_index <= 4977)) || ((pixel_index >= 4980) && (pixel_index <= 4981)) || ((pixel_index >= 5024) && (pixel_index <= 5026)) || ((pixel_index >= 5034) && (pixel_index <= 5035)) || ((pixel_index >= 5044) && (pixel_index <= 5045)) || ((pixel_index >= 5054) && (pixel_index <= 5055)) || ((pixel_index >= 5062) && (pixel_index <= 5063)) || ((pixel_index >= 5066) && (pixel_index <= 5067)) || ((pixel_index >= 5076) && (pixel_index <= 5077)) || ((pixel_index >= 5121) && (pixel_index <= 5123)) || ((pixel_index >= 5130) && (pixel_index <= 5131)) || ((pixel_index >= 5140) && (pixel_index <= 5141)) || ((pixel_index >= 5150) && (pixel_index <= 5151)) || ((pixel_index >= 5158) && (pixel_index <= 5159)) || ((pixel_index >= 5162) && (pixel_index <= 5163)) || ((pixel_index >= 5172) && (pixel_index <= 5173)) || ((pixel_index >= 5205) && (pixel_index <= 5220)) || ((pixel_index >= 5226) && (pixel_index <= 5227)) || ((pixel_index >= 5236) && (pixel_index <= 5241)) || ((pixel_index >= 5248) && (pixel_index <= 5249)) || ((pixel_index >= 5252) && (pixel_index <= 5253)) || ((pixel_index >= 5258) && (pixel_index <= 5263)) || ((pixel_index >= 5268) && (pixel_index <= 5269)) || ((pixel_index >= 5301) && (pixel_index <= 5316)) || ((pixel_index >= 5322) && (pixel_index <= 5323)) || ((pixel_index >= 5332) && (pixel_index <= 5337)) || ((pixel_index >= 5344) && (pixel_index <= 5345)) || ((pixel_index >= 5348) && (pixel_index <= 5349)) || ((pixel_index >= 5354) && (pixel_index <= 5359)) || ((pixel_index >= 5364) && (pixel_index <= 5365)) || ((pixel_index >= 5409) && (pixel_index <= 5411)) || ((pixel_index >= 5418) && (pixel_index <= 5419)) || ((pixel_index >= 5428) && (pixel_index <= 5429)) || ((pixel_index >= 5440) && (pixel_index <= 5441)) || ((pixel_index >= 5444) && (pixel_index <= 5445)) || ((pixel_index >= 5450) && (pixel_index <= 5451)) || ((pixel_index >= 5460) && (pixel_index <= 5461)) || ((pixel_index >= 5504) && (pixel_index <= 5506)) || ((pixel_index >= 5514) && (pixel_index <= 5515)) || ((pixel_index >= 5524) && (pixel_index <= 5525)) || ((pixel_index >= 5536) && (pixel_index <= 5537)) || ((pixel_index >= 5540) && (pixel_index <= 5541)) || ((pixel_index >= 5546) && (pixel_index <= 5547)) || ((pixel_index >= 5556) && (pixel_index <= 5557)) || ((pixel_index >= 5599) && (pixel_index <= 5601)) || ((pixel_index >= 5610) && (pixel_index <= 5617)) || ((pixel_index >= 5620) && (pixel_index <= 5627)) || ((pixel_index >= 5634) && (pixel_index <= 5635)) || ((pixel_index >= 5642) && (pixel_index <= 5649)) || ((pixel_index >= 5652) && (pixel_index <= 5659)) || ((pixel_index >= 5695) && (pixel_index <= 5696)) || ((pixel_index >= 5706) && (pixel_index <= 5713)) || ((pixel_index >= 5716) && (pixel_index <= 5723)) || ((pixel_index >= 5730) && (pixel_index <= 5731)) || ((pixel_index >= 5738) && (pixel_index <= 5745)) || (pixel_index >= 5748) && (pixel_index <= 5755)) oled_data = 16'b1111111111111111;
            else oled_data = 16'b0000000001000100;
        end
    end

endmodule

module gameoverbase_data(input [12:0] pixel_index, output reg [15:0] oled_data);
    wire [6:0] x = pixel_index % 96;
    wire [6:0] y = pixel_index / 96;
   
    always @ (*) begin
        if (((pixel_index >= 1159) && (pixel_index <= 1162)) || ((pixel_index >= 1169) && (pixel_index <= 1172)) || ((pixel_index >= 1177) && (pixel_index <= 1178)) || ((pixel_index >= 1185) && (pixel_index <= 1186)) || ((pixel_index >= 1189) && (pixel_index <= 1196)) || ((pixel_index >= 1205) && (pixel_index <= 1208)) || ((pixel_index >= 1213) && (pixel_index <= 1214)) || ((pixel_index >= 1221) && (pixel_index <= 1222)) || ((pixel_index >= 1225) && (pixel_index <= 1232)) || ((pixel_index >= 1235) && (pixel_index <= 1240)) || ((pixel_index >= 1255) && (pixel_index <= 1258)) || ((pixel_index >= 1265) && (pixel_index <= 1268)) || ((pixel_index >= 1273) && (pixel_index <= 1274)) || ((pixel_index >= 1281) && (pixel_index <= 1282)) || ((pixel_index >= 1285) && (pixel_index <= 1292)) || ((pixel_index >= 1301) && (pixel_index <= 1304)) || ((pixel_index >= 1309) && (pixel_index <= 1310)) || ((pixel_index >= 1317) && (pixel_index <= 1318)) || ((pixel_index >= 1321) && (pixel_index <= 1328)) || ((pixel_index >= 1331) && (pixel_index <= 1336)) || ((pixel_index >= 1349) && (pixel_index <= 1350)) || ((pixel_index >= 1359) && (pixel_index <= 1360)) || ((pixel_index >= 1365) && (pixel_index <= 1366)) || ((pixel_index >= 1369) && (pixel_index <= 1372)) || ((pixel_index >= 1375) && (pixel_index <= 1378)) || ((pixel_index >= 1381) && (pixel_index <= 1382)) || ((pixel_index >= 1395) && (pixel_index <= 1396)) || ((pixel_index >= 1401) && (pixel_index <= 1402)) || ((pixel_index >= 1405) && (pixel_index <= 1406)) || ((pixel_index >= 1413) && (pixel_index <= 1414)) || ((pixel_index >= 1417) && (pixel_index <= 1418)) || ((pixel_index >= 1427) && (pixel_index <= 1428)) || ((pixel_index >= 1433) && (pixel_index <= 1434)) || ((pixel_index >= 1445) && (pixel_index <= 1446)) || ((pixel_index >= 1455) && (pixel_index <= 1456)) || ((pixel_index >= 1461) && (pixel_index <= 1462)) || ((pixel_index >= 1465) && (pixel_index <= 1468)) || ((pixel_index >= 1471) && (pixel_index <= 1474)) || ((pixel_index >= 1477) && (pixel_index <= 1478)) || ((pixel_index >= 1491) && (pixel_index <= 1492)) || ((pixel_index >= 1497) && (pixel_index <= 1498)) || ((pixel_index >= 1501) && (pixel_index <= 1502)) || ((pixel_index >= 1509) && (pixel_index <= 1510)) || ((pixel_index >= 1513) && (pixel_index <= 1514)) || ((pixel_index >= 1523) && (pixel_index <= 1524)) || ((pixel_index >= 1529) && (pixel_index <= 1530)) || ((pixel_index >= 1541) && (pixel_index <= 1542)) || ((pixel_index >= 1545) && (pixel_index <= 1548)) || ((pixel_index >= 1551) && (pixel_index <= 1558)) || ((pixel_index >= 1561) && (pixel_index <= 1562)) || ((pixel_index >= 1565) && (pixel_index <= 1566)) || ((pixel_index >= 1569) && (pixel_index <= 1570)) || ((pixel_index >= 1573) && (pixel_index <= 1578)) || ((pixel_index >= 1587) && (pixel_index <= 1588)) || ((pixel_index >= 1593) && (pixel_index <= 1594)) || ((pixel_index >= 1599) && (pixel_index <= 1600)) || ((pixel_index >= 1603) && (pixel_index <= 1604)) || ((pixel_index >= 1609) && (pixel_index <= 1614)) || ((pixel_index >= 1619) && (pixel_index <= 1624)) || ((pixel_index >= 1637) && (pixel_index <= 1638)) || ((pixel_index >= 1641) && (pixel_index <= 1644)) || ((pixel_index >= 1647) && (pixel_index <= 1654)) || ((pixel_index >= 1657) && (pixel_index <= 1658)) || ((pixel_index >= 1661) && (pixel_index <= 1662)) || ((pixel_index >= 1665) && (pixel_index <= 1666)) || ((pixel_index >= 1669) && (pixel_index <= 1674)) || ((pixel_index >= 1683) && (pixel_index <= 1684)) || ((pixel_index >= 1689) && (pixel_index <= 1690)) || ((pixel_index >= 1695) && (pixel_index <= 1696)) || ((pixel_index >= 1699) && (pixel_index <= 1700)) || ((pixel_index >= 1705) && (pixel_index <= 1710)) || ((pixel_index >= 1715) && (pixel_index <= 1720)) || ((pixel_index >= 1733) && (pixel_index <= 1734)) || ((pixel_index >= 1739) && (pixel_index <= 1740)) || ((pixel_index >= 1743) && (pixel_index <= 1744)) || ((pixel_index >= 1749) && (pixel_index <= 1750)) || ((pixel_index >= 1753) && (pixel_index <= 1754)) || ((pixel_index >= 1761) && (pixel_index <= 1762)) || ((pixel_index >= 1765) && (pixel_index <= 1766)) || ((pixel_index >= 1779) && (pixel_index <= 1780)) || ((pixel_index >= 1785) && (pixel_index <= 1786)) || ((pixel_index >= 1791) && (pixel_index <= 1792)) || ((pixel_index >= 1795) && (pixel_index <= 1796)) || ((pixel_index >= 1801) && (pixel_index <= 1802)) || ((pixel_index >= 1811) && (pixel_index <= 1812)) || ((pixel_index >= 1815) && (pixel_index <= 1816)) || ((pixel_index >= 1829) && (pixel_index <= 1830)) || ((pixel_index >= 1835) && (pixel_index <= 1836)) || ((pixel_index >= 1839) && (pixel_index <= 1840)) || ((pixel_index >= 1845) && (pixel_index <= 1846)) || ((pixel_index >= 1849) && (pixel_index <= 1850)) || ((pixel_index >= 1857) && (pixel_index <= 1858)) || ((pixel_index >= 1861) && (pixel_index <= 1862)) || ((pixel_index >= 1875) && (pixel_index <= 1876)) || ((pixel_index >= 1881) && (pixel_index <= 1882)) || ((pixel_index >= 1887) && (pixel_index <= 1888)) || ((pixel_index >= 1891) && (pixel_index <= 1892)) || ((pixel_index >= 1897) && (pixel_index <= 1898)) || ((pixel_index >= 1907) && (pixel_index <= 1908)) || ((pixel_index >= 1911) && (pixel_index <= 1912)) || ((pixel_index >= 1927) && (pixel_index <= 1930)) || ((pixel_index >= 1935) && (pixel_index <= 1936)) || ((pixel_index >= 1941) && (pixel_index <= 1942)) || ((pixel_index >= 1945) && (pixel_index <= 1946)) || ((pixel_index >= 1953) && (pixel_index <= 1954)) || ((pixel_index >= 1957) && (pixel_index <= 1964)) || ((pixel_index >= 1973) && (pixel_index <= 1976)) || ((pixel_index >= 1985) && (pixel_index <= 1986)) || ((pixel_index >= 1993) && (pixel_index <= 2000)) || ((pixel_index >= 2003) && (pixel_index <= 2004)) || ((pixel_index >= 2009) && (pixel_index <= 2010)) || ((pixel_index >= 2023) && (pixel_index <= 2026)) || ((pixel_index >= 2031) && (pixel_index <= 2032)) || ((pixel_index >= 2037) && (pixel_index <= 2038)) || ((pixel_index >= 2041) && (pixel_index <= 2042)) || ((pixel_index >= 2049) && (pixel_index <= 2050)) || ((pixel_index >= 2053) && (pixel_index <= 2060)) || ((pixel_index >= 2069) && (pixel_index <= 2072)) || ((pixel_index >= 2081) && (pixel_index <= 2082)) || ((pixel_index >= 2089) && (pixel_index <= 2096)) || ((pixel_index >= 2099) && (pixel_index <= 2100)) || ((pixel_index >= 2105) && (pixel_index <= 2106)) || ((pixel_index >= 2626) && (pixel_index <= 2628)) || ((pixel_index >= 2638) && (pixel_index <= 2640)) || ((pixel_index >= 2644) && (pixel_index <= 2652)) || ((pixel_index >= 2656) && (pixel_index <= 2658)) || ((pixel_index >= 2665) && (pixel_index <= 2667)) || ((pixel_index >= 2674) && (pixel_index <= 2682)) || ((pixel_index >= 2722) && (pixel_index <= 2724)) || ((pixel_index >= 2734) && (pixel_index <= 2736)) || ((pixel_index >= 2740) && (pixel_index <= 2748)) || ((pixel_index >= 2752) && (pixel_index <= 2754)) || ((pixel_index >= 2761) && (pixel_index <= 2763)) || ((pixel_index >= 2770) && (pixel_index <= 2778)) || ((pixel_index >= 2818) && (pixel_index <= 2820)) || ((pixel_index >= 2830) && (pixel_index <= 2832)) || ((pixel_index >= 2836) && (pixel_index <= 2844)) || ((pixel_index >= 2848) && (pixel_index <= 2850)) || ((pixel_index >= 2857) && (pixel_index <= 2859)) || ((pixel_index >= 2866) && (pixel_index <= 2874)) || ((pixel_index >= 2914) && (pixel_index <= 2916)) || ((pixel_index >= 2926) && (pixel_index <= 2928)) || ((pixel_index >= 2935) && (pixel_index <= 2937)) || ((pixel_index >= 2944) && (pixel_index <= 2949)) || ((pixel_index >= 2953) && (pixel_index <= 2955)) || ((pixel_index >= 2959) && (pixel_index <= 2961)) || ((pixel_index >= 3010) && (pixel_index <= 3012)) || ((pixel_index >= 3022) && (pixel_index <= 3024)) || ((pixel_index >= 3031) && (pixel_index <= 3033)) || ((pixel_index >= 3040) && (pixel_index <= 3045)) || ((pixel_index >= 3049) && (pixel_index <= 3051)) || ((pixel_index >= 3055) && (pixel_index <= 3057)) || ((pixel_index >= 3106) && (pixel_index <= 3108)) || ((pixel_index >= 3118) && (pixel_index <= 3120)) || ((pixel_index >= 3127) && (pixel_index <= 3129)) || ((pixel_index >= 3136) && (pixel_index <= 3141)) || ((pixel_index >= 3145) && (pixel_index <= 3147)) || ((pixel_index >= 3151) && (pixel_index <= 3153)) || ((pixel_index >= 3202) && (pixel_index <= 3204)) || ((pixel_index >= 3208) && (pixel_index <= 3210)) || ((pixel_index >= 3214) && (pixel_index <= 3216)) || ((pixel_index >= 3223) && (pixel_index <= 3225)) || ((pixel_index >= 3232) && (pixel_index <= 3234)) || ((pixel_index >= 3238) && (pixel_index <= 3243)) || ((pixel_index >= 3250) && (pixel_index <= 3255)) || ((pixel_index >= 3298) && (pixel_index <= 3300)) || ((pixel_index >= 3304) && (pixel_index <= 3306)) || ((pixel_index >= 3310) && (pixel_index <= 3312)) || ((pixel_index >= 3319) && (pixel_index <= 3321)) || ((pixel_index >= 3328) && (pixel_index <= 3330)) || ((pixel_index >= 3334) && (pixel_index <= 3339)) || ((pixel_index >= 3346) && (pixel_index <= 3351)) || ((pixel_index >= 3394) && (pixel_index <= 3396)) || ((pixel_index >= 3400) && (pixel_index <= 3402)) || ((pixel_index >= 3406) && (pixel_index <= 3408)) || ((pixel_index >= 3415) && (pixel_index <= 3417)) || ((pixel_index >= 3424) && (pixel_index <= 3426)) || ((pixel_index >= 3430) && (pixel_index <= 3435)) || ((pixel_index >= 3442) && (pixel_index <= 3447)) || ((pixel_index >= 3490) && (pixel_index <= 3495)) || ((pixel_index >= 3499) && (pixel_index <= 3504)) || ((pixel_index >= 3511) && (pixel_index <= 3513)) || ((pixel_index >= 3520) && (pixel_index <= 3522)) || ((pixel_index >= 3529) && (pixel_index <= 3531)) || ((pixel_index >= 3544) && (pixel_index <= 3546)) || ((pixel_index >= 3586) && (pixel_index <= 3591)) || ((pixel_index >= 3595) && (pixel_index <= 3600)) || ((pixel_index >= 3607) && (pixel_index <= 3609)) || ((pixel_index >= 3616) && (pixel_index <= 3618)) || ((pixel_index >= 3625) && (pixel_index <= 3627)) || ((pixel_index >= 3640) && (pixel_index <= 3642)) || ((pixel_index >= 3682) && (pixel_index <= 3687)) || ((pixel_index >= 3691) && (pixel_index <= 3696)) || ((pixel_index >= 3703) && (pixel_index <= 3705)) || ((pixel_index >= 3712) && (pixel_index <= 3714)) || ((pixel_index >= 3721) && (pixel_index <= 3723)) || ((pixel_index >= 3736) && (pixel_index <= 3738)) || ((pixel_index >= 3778) && (pixel_index <= 3780)) || ((pixel_index >= 3790) && (pixel_index <= 3792)) || ((pixel_index >= 3796) && (pixel_index <= 3804)) || ((pixel_index >= 3808) && (pixel_index <= 3810)) || ((pixel_index >= 3817) && (pixel_index <= 3819)) || ((pixel_index >= 3823) && (pixel_index <= 3831)) || ((pixel_index >= 3874) && (pixel_index <= 3876)) || ((pixel_index >= 3886) && (pixel_index <= 3888)) || ((pixel_index >= 3892) && (pixel_index <= 3900)) || ((pixel_index >= 3904) && (pixel_index <= 3906)) || ((pixel_index >= 3913) && (pixel_index <= 3915)) || ((pixel_index >= 3919) && (pixel_index <= 3927)) || ((pixel_index >= 3970) && (pixel_index <= 3972)) || ((pixel_index >= 3982) && (pixel_index <= 3984)) || ((pixel_index >= 3988) && (pixel_index <= 3996)) || ((pixel_index >= 4000) && (pixel_index <= 4002)) || ((pixel_index >= 4009) && (pixel_index <= 4011)) || (pixel_index >= 4015) && (pixel_index <= 4023)) oled_data = 16'b1111111111111111;
        else if (x <= 30 && y >= 26 && y <= 51) oled_data = 0;
        else oled_data = 16'b0000000001000100;
    end

endmodule

module gameoverresult_data(input sw, input [12:0] pixel_index, output reg [15:0] oled_data);
    wire [6:0] x = pixel_index % 96;
    wire [6:0] y = pixel_index / 96;
    
    always @ (*) begin
        if (x >= 31 && y <= 25 && y >= 52) oled_data = 0;
        if (sw == 0) begin // cross
            if (((pixel_index >= 2502) && (pixel_index <= 2504)) || ((pixel_index >= 2523) && (pixel_index <= 2525)) || ((pixel_index >= 2597) && (pixel_index <= 2601)) || pixel_index == 2618 || ((pixel_index >= 2620) && (pixel_index <= 2622)) || ((pixel_index >= 2693) && (pixel_index <= 2694)) || ((pixel_index >= 2696) && (pixel_index <= 2698)) || ((pixel_index >= 2713) && (pixel_index <= 2718)) || ((pixel_index >= 2789) && (pixel_index <= 2792)) || ((pixel_index >= 2794) && (pixel_index <= 2795)) || ((pixel_index >= 2808) && (pixel_index <= 2809)) || pixel_index == 2811 || pixel_index == 2813 || pixel_index == 2886 || ((pixel_index >= 2888) && (pixel_index <= 2892)) || ((pixel_index >= 2903) && (pixel_index <= 2909)) || ((pixel_index >= 2983) && (pixel_index <= 2986)) || ((pixel_index >= 2988) && (pixel_index <= 2989)) || ((pixel_index >= 2998) && (pixel_index <= 3000)) || ((pixel_index >= 3002) && (pixel_index <= 3004)) || pixel_index == 3080 || ((pixel_index >= 3082) && (pixel_index <= 3086)) || pixel_index == 3093 || ((pixel_index >= 3095) && (pixel_index <= 3098)) || ((pixel_index >= 3177) && (pixel_index <= 3179)) || ((pixel_index >= 3181) && (pixel_index <= 3183)) || ((pixel_index >= 3188) && (pixel_index <= 3191)) || ((pixel_index >= 3193) && (pixel_index <= 3194)) || ((pixel_index >= 3274) && (pixel_index <= 3277)) || ((pixel_index >= 3279) && (pixel_index <= 3280)) || ((pixel_index >= 3283) && (pixel_index <= 3285)) || ((pixel_index >= 3287) && (pixel_index <= 3289)) || ((pixel_index >= 3371) && (pixel_index <= 3372)) || ((pixel_index >= 3374) && (pixel_index <= 3378)) || ((pixel_index >= 3380) && (pixel_index <= 3383)) || ((pixel_index >= 3469) && (pixel_index <= 3470)) || ((pixel_index >= 3472) && (pixel_index <= 3476)) || ((pixel_index >= 3478) && (pixel_index <= 3479)) || ((pixel_index >= 3565) && (pixel_index <= 3568)) || ((pixel_index >= 3570) && (pixel_index <= 3574)) || ((pixel_index >= 3662) && (pixel_index <= 3666)) || pixel_index == 3668 || pixel_index == 3758 || pixel_index == 3760 || ((pixel_index >= 3762) && (pixel_index <= 3763)) || pixel_index == 3765 || ((pixel_index >= 3854) && (pixel_index <= 3859)) || ((pixel_index >= 3861) && (pixel_index <= 3862)) || ((pixel_index >= 3948) && (pixel_index <= 3951)) || ((pixel_index >= 3953) && (pixel_index <= 3959)) || ((pixel_index >= 4043) && (pixel_index <= 4045)) || ((pixel_index >= 4047) && (pixel_index <= 4049)) || ((pixel_index >= 4051) && (pixel_index <= 4052)) || ((pixel_index >= 4054) && (pixel_index <= 4056)) || ((pixel_index >= 4138) && (pixel_index <= 4140)) || ((pixel_index >= 4142) && (pixel_index <= 4144)) || ((pixel_index >= 4147) && (pixel_index <= 4150)) || ((pixel_index >= 4152) && (pixel_index <= 4153)) || ((pixel_index >= 4233) && (pixel_index <= 4239)) || ((pixel_index >= 4244) && (pixel_index <= 4250)) || ((pixel_index >= 4328) && (pixel_index <= 4330)) || ((pixel_index >= 4332) && (pixel_index <= 4333)) || pixel_index == 4341 || ((pixel_index >= 4343) && (pixel_index <= 4344)) || ((pixel_index >= 4346) && (pixel_index <= 4347)) || ((pixel_index >= 4423) && (pixel_index <= 4429)) || ((pixel_index >= 4438) && (pixel_index <= 4444)) || pixel_index == 4518 || ((pixel_index >= 4520) && (pixel_index <= 4521)) || pixel_index == 4523 || pixel_index == 4536 || ((pixel_index >= 4538) && (pixel_index <= 4541)) || ((pixel_index >= 4613) && (pixel_index <= 4617)) || pixel_index == 4619 || pixel_index == 4632 || pixel_index == 4634 || ((pixel_index >= 4636) && (pixel_index <= 4638)) || ((pixel_index >= 4709) && (pixel_index <= 4710)) || pixel_index == 4712 || pixel_index == 4714 || ((pixel_index >= 4729) && (pixel_index <= 4732)) || pixel_index == 4734 || ((pixel_index >= 4805) && (pixel_index <= 4809)) || ((pixel_index >= 4827) && (pixel_index <= 4830)) || ((pixel_index >= 4903) && (pixel_index <= 4904)) || (pixel_index >= 4923) && (pixel_index <= 4924) || pixel_index == 2619 || pixel_index == 2695 || pixel_index == 2793 || pixel_index == 2810 || pixel_index == 2812 || pixel_index == 2814 || pixel_index == 2887 || pixel_index == 2987 || pixel_index == 3001 || pixel_index == 3081 || pixel_index == 3094 || pixel_index == 3099 || pixel_index == 3180 || pixel_index == 3192 || pixel_index == 3278 || pixel_index == 3286 || pixel_index == 3379 || pixel_index == 3468 || pixel_index == 3471 || pixel_index == 3477 || pixel_index == 3569 || pixel_index == 3667 || pixel_index == 3669 || pixel_index == 3759 || pixel_index == 3761 || pixel_index == 3853 || pixel_index == 3860 || pixel_index == 3952 || pixel_index == 4046 || pixel_index == 4050 || pixel_index == 4053 || pixel_index == 4141 || pixel_index == 4151 || pixel_index == 4331 || pixel_index == 4334 || pixel_index == 4342 || pixel_index == 4345 || pixel_index == 4519 || pixel_index == 4522 || pixel_index == 4524 || pixel_index == 4535 || pixel_index == 4537 || pixel_index == 4635 || pixel_index == 4711 || pixel_index == 4713 || pixel_index == 4733 || pixel_index == 4826 || pixel_index == 4902 || pixel_index == 4925 || pixel_index == 3373 || pixel_index == 3384 || pixel_index == 3764 || pixel_index == 4618 || pixel_index == 4633) oled_data = 16'b0001011101111111;
            else oled_data = 16'b0000000001000100;
        end
        if (sw == 1) begin // circle
            if (pixel_index == 2509 || ((pixel_index >= 2511) && (pixel_index <= 2512)) || ((pixel_index >= 2514) && (pixel_index <= 2515)) || ((pixel_index >= 2517) && (pixel_index <= 2518)) || pixel_index == 2604 || pixel_index == 2606 || pixel_index == 2609 || ((pixel_index >= 2611) && (pixel_index <= 2612)) || pixel_index == 2614 || pixel_index == 2616 || ((pixel_index >= 2699) && (pixel_index <= 2701)) || pixel_index == 2703 || ((pixel_index >= 2705) && (pixel_index <= 2706)) || pixel_index == 2708 || ((pixel_index >= 2710) && (pixel_index <= 2711)) || pixel_index == 2713 || ((pixel_index >= 2793) && (pixel_index <= 2794)) || pixel_index == 2796 || ((pixel_index >= 2798) && (pixel_index <= 2800)) || pixel_index == 2802 || ((pixel_index >= 2804) && (pixel_index <= 2805)) || pixel_index == 2807 || pixel_index == 2809 || pixel_index == 2889 || pixel_index == 2891 || ((pixel_index >= 2893) && (pixel_index <= 2894)) || pixel_index == 2902 || pixel_index == 2904 || ((pixel_index >= 2906) && (pixel_index <= 2907)) || pixel_index == 2985 || ((pixel_index >= 2987) && (pixel_index <= 2988)) || ((pixel_index >= 2999) && (pixel_index <= 3001)) || pixel_index == 3003 || pixel_index == 3079 || pixel_index == 3081 || pixel_index == 3084 || pixel_index == 3095 || ((pixel_index >= 3097) && (pixel_index <= 3098)) || pixel_index == 3100 || ((pixel_index >= 3174) && (pixel_index <= 3175)) || pixel_index == 3177 || pixel_index == 3179 || pixel_index == 3193 || ((pixel_index >= 3195) && (pixel_index <= 3197)) || ((pixel_index >= 3272) && (pixel_index <= 3274)) || pixel_index == 3289 || pixel_index == 3293 || pixel_index == 3365 || pixel_index == 3367 || pixel_index == 3369 || pixel_index == 3386 || pixel_index == 3388 || pixel_index == 3390 || ((pixel_index >= 3462) && (pixel_index <= 3464)) || ((pixel_index >= 3483) && (pixel_index <= 3484)) || pixel_index == 3557 || ((pixel_index >= 3581) && (pixel_index <= 3582)) || pixel_index == 3654 || pixel_index == 3656 || pixel_index == 3676 || pixel_index == 3678 || ((pixel_index >= 3749) && (pixel_index <= 3751)) || pixel_index == 3771 || pixel_index == 3773 || pixel_index == 3846 || pixel_index == 3848 || ((pixel_index >= 3868) && (pixel_index <= 3870)) || ((pixel_index >= 3942) && (pixel_index <= 3943)) || pixel_index == 3945 || pixel_index == 3963 || pixel_index == 4037 || pixel_index == 4039 || pixel_index == 4058 || ((pixel_index >= 4060) && (pixel_index <= 4061)) || pixel_index == 4133 || pixel_index == 4135 || pixel_index == 4137 || pixel_index == 4154 || ((pixel_index >= 4157) && (pixel_index <= 4158)) || pixel_index == 4230 || pixel_index == 4232 || pixel_index == 4234 || pixel_index == 4249 || ((pixel_index >= 4251) && (pixel_index <= 4252)) || pixel_index == 4327 || pixel_index == 4329 || pixel_index == 4331 || pixel_index == 4344 || ((pixel_index >= 4348) && (pixel_index <= 4349)) || pixel_index == 4423 || ((pixel_index >= 4426) && (pixel_index <= 4429)) || pixel_index == 4439 || ((pixel_index >= 4441) && (pixel_index <= 4443)) || pixel_index == 4521 || pixel_index == 4523 || pixel_index == 4527 || ((pixel_index >= 4533) && (pixel_index <= 4534)) || pixel_index == 4537 || pixel_index == 4539 || pixel_index == 4616 || ((pixel_index >= 4618) && (pixel_index <= 4619)) || pixel_index == 4621 || pixel_index == 4623 || pixel_index == 4625 || ((pixel_index >= 4627) && (pixel_index <= 4628)) || ((pixel_index >= 4630) && (pixel_index <= 4631)) || pixel_index == 4633 || pixel_index == 4635 || ((pixel_index >= 4715) && (pixel_index <= 4716)) || ((pixel_index >= 4718) && (pixel_index <= 4719)) || pixel_index == 4721 || pixel_index == 4725 || ((pixel_index >= 4727) && (pixel_index <= 4728)) || pixel_index == 4812 || pixel_index == 4816 || ((pixel_index >= 4818) && (pixel_index <= 4820)) || pixel_index == 4822 || pixel_index == 4824 || pixel_index == 4910 || pixel_index == 4912 || pixel_index == 4915 || pixel_index == 4918 || pixel_index == 2510 || pixel_index == 2513 || pixel_index == 2516 || pixel_index == 2603 || pixel_index == 2605 || pixel_index == 2607 || pixel_index == 2610 || pixel_index == 2615 || pixel_index == 2698 || pixel_index == 2704 || pixel_index == 2709 || pixel_index == 2712 || pixel_index == 2792 || pixel_index == 2795 || pixel_index == 2797 || pixel_index == 2801 || pixel_index == 2803 || pixel_index == 2806 || ((pixel_index >= 2810) && (pixel_index <= 2811)) || pixel_index == 2888 || pixel_index == 2890 || pixel_index == 2895 || pixel_index == 2900 || pixel_index == 2903 || pixel_index == 2905 || pixel_index == 2983 || pixel_index == 2986 || pixel_index == 2989 || pixel_index == 2998 || pixel_index == 3004 || pixel_index == 3078 || pixel_index == 3080 || pixel_index == 3083 || pixel_index == 3099 || pixel_index == 3101 || pixel_index == 3178 || pixel_index == 3192 || pixel_index == 3194 || pixel_index == 3269 || pixel_index == 3271 || pixel_index == 3290 || pixel_index == 3292 || pixel_index == 3366 || pixel_index == 3368 || pixel_index == 3387 || pixel_index == 3389 || pixel_index == 3461 || pixel_index == 3465 || pixel_index == 3482 || pixel_index == 3486 || pixel_index == 3558 || pixel_index == 3560 || pixel_index == 3580 || pixel_index == 3653 || pixel_index == 3655 || pixel_index == 3675 || pixel_index == 3677 || pixel_index == 3752 || pixel_index == 3772 || pixel_index == 3845 || pixel_index == 3867 || pixel_index == 3941 || pixel_index == 3944 || pixel_index == 3962 || pixel_index == 3964 || pixel_index == 3966 || pixel_index == 4038 || pixel_index == 4041 || pixel_index == 4059 || pixel_index == 4062 || pixel_index == 4134 || pixel_index == 4136 || pixel_index == 4138 || pixel_index == 4153 || pixel_index == 4156 || pixel_index == 4231 || pixel_index == 4235 || pixel_index == 4248 || pixel_index == 4250 || pixel_index == 4253 || pixel_index == 4326 || pixel_index == 4328 || pixel_index == 4330 || pixel_index == 4332 || pixel_index == 4345 || pixel_index == 4347 || pixel_index == 4425 || pixel_index == 4438 || pixel_index == 4440 || pixel_index == 4520 || pixel_index == 4524 || pixel_index == 4526 || pixel_index == 4532 || pixel_index == 4535 || pixel_index == 4538 || pixel_index == 4617 || pixel_index == 4620 || pixel_index == 4622 || pixel_index == 4624 || pixel_index == 4626 || pixel_index == 4632 || pixel_index == 4634 || pixel_index == 4714 || pixel_index == 4717 || pixel_index == 4720 || pixel_index == 4722 || pixel_index == 4724 || pixel_index == 4726 || pixel_index == 4814 || pixel_index == 4817 || pixel_index == 4821 || pixel_index == 4909 || pixel_index == 4911 || pixel_index == 4914 || pixel_index == 4916 || pixel_index == 2608 || pixel_index == 2901 || pixel_index == 2984 || pixel_index == 3082 || pixel_index == 3270 || pixel_index == 3291 || pixel_index == 3485 || pixel_index == 3559 || pixel_index == 3579 || pixel_index == 3965 || pixel_index == 4040 || pixel_index == 4155 || pixel_index == 4233 || pixel_index == 4343 || pixel_index == 4346 || pixel_index == 4424 || pixel_index == 4525 || pixel_index == 4536 || pixel_index == 4723 || pixel_index == 4813 || pixel_index == 4815 || pixel_index == 4913 || pixel_index == 4917 || pixel_index == 2613 || pixel_index == 2702 || pixel_index == 2707 || pixel_index == 2808 || pixel_index == 2892 || pixel_index == 3002 || pixel_index == 3096 || pixel_index == 3176 || pixel_index == 3294 || pixel_index == 3774 || pixel_index == 3847 || pixel_index == 4444 || pixel_index == 4522 || pixel_index == 4629 || pixel_index == 4729 || pixel_index == 4811 || pixel_index == 4823) oled_data = 16'b1111100001011010;
            else oled_data = 16'b0000000001000100;
        end
    end

endmodule

module x_win_anim(input frame_rate, input start, input [12:0] pixel_index, output reg done, output reg [15:0] oled_data);
    reg [15:0] frame_count = 0;
    
    always @ (posedge frame_rate) begin
        if (start) frame_count <= (frame_count == 31) ? 31 : frame_count + 1;
        else frame_count <= 0;
    end
   
    // animation for X win (1v1 mode) or player win (AI mode)
    // Reimu throwing apple up
    always @ (*) begin
        if (frame_count <= 30) done = 0;
        if (frame_count == 0) oled_data = 0;
        else if (frame_count == 1) begin
            if (((pixel_index >= 5) && (pixel_index <= 54)) || ((pixel_index >= 61) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 150)) || ((pixel_index >= 158) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 245)) || ((pixel_index >= 255) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 342)) || ((pixel_index >= 352) && (pixel_index <= 377)) || ((pixel_index >= 389) && (pixel_index <= 438)) || ((pixel_index >= 449) && (pixel_index <= 451)) || ((pixel_index >= 453) && (pixel_index <= 473)) || ((pixel_index >= 485) && (pixel_index <= 534)) || ((pixel_index >= 552) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 631)) || ((pixel_index >= 649) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 726)) || ((pixel_index >= 746) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 820)) || ((pixel_index >= 842) && (pixel_index <= 857)) || ((pixel_index >= 869) && (pixel_index <= 914)) || ((pixel_index >= 939) && (pixel_index <= 953)) || ((pixel_index >= 965) && (pixel_index <= 1009)) || ((pixel_index >= 1035) && (pixel_index <= 1049)) || ((pixel_index >= 1061) && (pixel_index <= 1104)) || ((pixel_index >= 1131) && (pixel_index <= 1145)) || ((pixel_index >= 1157) && (pixel_index <= 1199)) || ((pixel_index >= 1228) && (pixel_index <= 1241)) || ((pixel_index >= 1253) && (pixel_index <= 1295)) || ((pixel_index >= 1324) && (pixel_index <= 1337)) || ((pixel_index >= 1349) && (pixel_index <= 1390)) || ((pixel_index >= 1421) && (pixel_index <= 1433)) || ((pixel_index >= 1445) && (pixel_index <= 1486)) || ((pixel_index >= 1517) && (pixel_index <= 1529)) || ((pixel_index >= 1541) && (pixel_index <= 1581)) || ((pixel_index >= 1613) && (pixel_index <= 1625)) || ((pixel_index >= 1637) && (pixel_index <= 1677)) || ((pixel_index >= 1710) && (pixel_index <= 1721)) || ((pixel_index >= 1733) && (pixel_index <= 1773)) || ((pixel_index >= 1806) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1869)) || ((pixel_index >= 1902) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 1965)) || ((pixel_index >= 1998) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2061)) || ((pixel_index >= 2095) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2157)) || ((pixel_index >= 2191) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2254)) || ((pixel_index >= 2287) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2351)) || ((pixel_index >= 2383) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2448)) || ((pixel_index >= 2479) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2546)) || ((pixel_index >= 2575) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2642)) || ((pixel_index >= 2671) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2737)) || ((pixel_index >= 2767) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2833)) || ((pixel_index >= 2863) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2930)) || ((pixel_index >= 2960) && (pixel_index <= 2969)) || ((pixel_index >= 2981) && (pixel_index <= 3027)) || ((pixel_index >= 3056) && (pixel_index <= 3065)) || ((pixel_index >= 3077) && (pixel_index <= 3124)) || ((pixel_index >= 3151) && (pixel_index <= 3161)) || ((pixel_index >= 3173) && (pixel_index <= 3220)) || ((pixel_index >= 3248) && (pixel_index <= 3257)) || ((pixel_index >= 3269) && (pixel_index <= 3317)) || ((pixel_index >= 3344) && (pixel_index <= 3353)) || ((pixel_index >= 3365) && (pixel_index <= 3413)) || ((pixel_index >= 3440) && (pixel_index <= 3449)) || ((pixel_index >= 3461) && (pixel_index <= 3492)) || ((pixel_index >= 3497) && (pixel_index <= 3509)) || ((pixel_index >= 3536) && (pixel_index <= 3545)) || ((pixel_index >= 3557) && (pixel_index <= 3586)) || ((pixel_index >= 3595) && (pixel_index <= 3605)) || ((pixel_index >= 3632) && (pixel_index <= 3641)) || ((pixel_index >= 3653) && (pixel_index <= 3680)) || ((pixel_index >= 3691) && (pixel_index <= 3701)) || ((pixel_index >= 3728) && (pixel_index <= 3737)) || ((pixel_index >= 3749) && (pixel_index <= 3775)) || ((pixel_index >= 3787) && (pixel_index <= 3798)) || ((pixel_index >= 3824) && (pixel_index <= 3833)) || ((pixel_index >= 3845) && (pixel_index <= 3871)) || ((pixel_index >= 3884) && (pixel_index <= 3894)) || ((pixel_index >= 3920) && (pixel_index <= 3929)) || ((pixel_index >= 3941) && (pixel_index <= 3967)) || ((pixel_index >= 3980) && (pixel_index <= 3990)) || pixel_index == 4012 || ((pixel_index >= 4016) && (pixel_index <= 4025)) || ((pixel_index >= 4037) && (pixel_index <= 4063)) || ((pixel_index >= 4076) && (pixel_index <= 4086)) || ((pixel_index >= 4108) && (pixel_index <= 4110)) || ((pixel_index >= 4112) && (pixel_index <= 4121)) || ((pixel_index >= 4133) && (pixel_index <= 4159)) || ((pixel_index >= 4172) && (pixel_index <= 4182)) || ((pixel_index >= 4203) && (pixel_index <= 4217)) || ((pixel_index >= 4229) && (pixel_index <= 4255)) || ((pixel_index >= 4268) && (pixel_index <= 4278)) || ((pixel_index >= 4299) && (pixel_index <= 4313)) || ((pixel_index >= 4325) && (pixel_index <= 4351)) || ((pixel_index >= 4365) && (pixel_index <= 4374)) || ((pixel_index >= 4395) && (pixel_index <= 4409)) || ((pixel_index >= 4421) && (pixel_index <= 4448)) || ((pixel_index >= 4462) && (pixel_index <= 4466)) || ((pixel_index >= 4468) && (pixel_index <= 4469)) || ((pixel_index >= 4491) && (pixel_index <= 4505)) || ((pixel_index >= 4517) && (pixel_index <= 4545)) || ((pixel_index >= 4559) && (pixel_index <= 4561)) || pixel_index == 4585 || ((pixel_index >= 4588) && (pixel_index <= 4601)) || ((pixel_index >= 4613) && (pixel_index <= 4641)) || ((pixel_index >= 4656) && (pixel_index <= 4657)) || ((pixel_index >= 4682) && (pixel_index <= 4697)) || ((pixel_index >= 4709) && (pixel_index <= 4739)) || ((pixel_index >= 4752) && (pixel_index <= 4753)) || ((pixel_index >= 4778) && (pixel_index <= 4793)) || ((pixel_index >= 4805) && (pixel_index <= 4837)) || pixel_index == 4849 || ((pixel_index >= 4874) && (pixel_index <= 4889)) || ((pixel_index >= 4901) && (pixel_index <= 4933)) || ((pixel_index >= 4970) && (pixel_index <= 4985)) || ((pixel_index >= 4997) && (pixel_index <= 5028)) || ((pixel_index >= 5066) && (pixel_index <= 5081)) || ((pixel_index >= 5093) && (pixel_index <= 5124)) || ((pixel_index >= 5163) && (pixel_index <= 5177)) || ((pixel_index >= 5189) && (pixel_index <= 5220)) || ((pixel_index >= 5259) && (pixel_index <= 5273)) || ((pixel_index >= 5285) && (pixel_index <= 5315)) || ((pixel_index >= 5355) && (pixel_index <= 5369)) || ((pixel_index >= 5381) && (pixel_index <= 5411)) || ((pixel_index >= 5451) && (pixel_index <= 5465)) || ((pixel_index >= 5477) && (pixel_index <= 5507)) || ((pixel_index >= 5547) && (pixel_index <= 5551)) || ((pixel_index >= 5553) && (pixel_index <= 5561)) || ((pixel_index >= 5573) && (pixel_index <= 5603)) || ((pixel_index >= 5644) && (pixel_index <= 5645)) || ((pixel_index >= 5649) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5699)) || ((pixel_index >= 5745) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5795)) || ((pixel_index >= 5838) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5891)) || ((pixel_index >= 5933) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 5986)) || pixel_index == 6005 || ((pixel_index >= 6029) && (pixel_index <= 6041)) || ((pixel_index >= 6053) && (pixel_index <= 6082)) || ((pixel_index >= 6101) && (pixel_index <= 6102)) || (pixel_index >= 6126) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 2) begin
            if (((pixel_index >= 5) && (pixel_index <= 55)) || ((pixel_index >= 65) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 150)) || ((pixel_index >= 162) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 247)) || ((pixel_index >= 259) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 343)) || ((pixel_index >= 355) && (pixel_index <= 356)) || ((pixel_index >= 359) && (pixel_index <= 377)) || ((pixel_index >= 389) && (pixel_index <= 439)) || ((pixel_index >= 457) && (pixel_index <= 473)) || ((pixel_index >= 485) && (pixel_index <= 536)) || ((pixel_index >= 554) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 630)) || ((pixel_index >= 651) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 724)) || ((pixel_index >= 748) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 818)) || ((pixel_index >= 844) && (pixel_index <= 857)) || ((pixel_index >= 869) && (pixel_index <= 913)) || ((pixel_index >= 941) && (pixel_index <= 953)) || ((pixel_index >= 965) && (pixel_index <= 1008)) || ((pixel_index >= 1037) && (pixel_index <= 1049)) || ((pixel_index >= 1061) && (pixel_index <= 1103)) || ((pixel_index >= 1133) && (pixel_index <= 1145)) || ((pixel_index >= 1157) && (pixel_index <= 1199)) || ((pixel_index >= 1230) && (pixel_index <= 1241)) || ((pixel_index >= 1253) && (pixel_index <= 1294)) || ((pixel_index >= 1326) && (pixel_index <= 1337)) || ((pixel_index >= 1349) && (pixel_index <= 1390)) || ((pixel_index >= 1423) && (pixel_index <= 1433)) || ((pixel_index >= 1445) && (pixel_index <= 1485)) || ((pixel_index >= 1519) && (pixel_index <= 1529)) || ((pixel_index >= 1541) && (pixel_index <= 1581)) || ((pixel_index >= 1615) && (pixel_index <= 1625)) || ((pixel_index >= 1637) && (pixel_index <= 1677)) || ((pixel_index >= 1712) && (pixel_index <= 1721)) || ((pixel_index >= 1733) && (pixel_index <= 1772)) || ((pixel_index >= 1808) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1869)) || ((pixel_index >= 1904) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 1965)) || ((pixel_index >= 2000) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2061)) || ((pixel_index >= 2096) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2157)) || ((pixel_index >= 2193) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2254)) || ((pixel_index >= 2289) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2351)) || ((pixel_index >= 2385) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2449)) || ((pixel_index >= 2481) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2546)) || ((pixel_index >= 2577) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2642)) || ((pixel_index >= 2673) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2737)) || ((pixel_index >= 2769) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2833)) || ((pixel_index >= 2865) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2930)) || ((pixel_index >= 2961) && (pixel_index <= 2969)) || ((pixel_index >= 2981) && (pixel_index <= 3027)) || ((pixel_index >= 3058) && (pixel_index <= 3065)) || ((pixel_index >= 3077) && (pixel_index <= 3124)) || ((pixel_index >= 3154) && (pixel_index <= 3161)) || ((pixel_index >= 3173) && (pixel_index <= 3220)) || ((pixel_index >= 3250) && (pixel_index <= 3257)) || ((pixel_index >= 3269) && (pixel_index <= 3317)) || ((pixel_index >= 3346) && (pixel_index <= 3353)) || ((pixel_index >= 3365) && (pixel_index <= 3397)) || ((pixel_index >= 3404) && (pixel_index <= 3413)) || ((pixel_index >= 3442) && (pixel_index <= 3449)) || ((pixel_index >= 3461) && (pixel_index <= 3490)) || ((pixel_index >= 3501) && (pixel_index <= 3509)) || ((pixel_index >= 3538) && (pixel_index <= 3545)) || ((pixel_index >= 3557) && (pixel_index <= 3585)) || ((pixel_index >= 3597) && (pixel_index <= 3605)) || ((pixel_index >= 3634) && (pixel_index <= 3641)) || ((pixel_index >= 3653) && (pixel_index <= 3681)) || ((pixel_index >= 3694) && (pixel_index <= 3702)) || ((pixel_index >= 3730) && (pixel_index <= 3737)) || ((pixel_index >= 3749) && (pixel_index <= 3777)) || ((pixel_index >= 3790) && (pixel_index <= 3798)) || ((pixel_index >= 3826) && (pixel_index <= 3833)) || ((pixel_index >= 3845) && (pixel_index <= 3872)) || ((pixel_index >= 3886) && (pixel_index <= 3894)) || pixel_index == 3917 || ((pixel_index >= 3922) && (pixel_index <= 3929)) || ((pixel_index >= 3941) && (pixel_index <= 3968)) || ((pixel_index >= 3982) && (pixel_index <= 3990)) || ((pixel_index >= 4018) && (pixel_index <= 4025)) || ((pixel_index >= 4037) && (pixel_index <= 4065)) || ((pixel_index >= 4078) && (pixel_index <= 4087)) || pixel_index == 4110 || pixel_index == 4112 || ((pixel_index >= 4114) && (pixel_index <= 4121)) || ((pixel_index >= 4133) && (pixel_index <= 4161)) || ((pixel_index >= 4174) && (pixel_index <= 4183)) || ((pixel_index >= 4206) && (pixel_index <= 4217)) || ((pixel_index >= 4229) && (pixel_index <= 4257)) || ((pixel_index >= 4271) && (pixel_index <= 4279)) || ((pixel_index >= 4301) && (pixel_index <= 4313)) || ((pixel_index >= 4325) && (pixel_index <= 4353)) || ((pixel_index >= 4368) && (pixel_index <= 4374)) || ((pixel_index >= 4397) && (pixel_index <= 4409)) || ((pixel_index >= 4421) && (pixel_index <= 4450)) || ((pixel_index >= 4465) && (pixel_index <= 4470)) || ((pixel_index >= 4493) && (pixel_index <= 4505)) || ((pixel_index >= 4517) && (pixel_index <= 4547)) || ((pixel_index >= 4564) && (pixel_index <= 4565)) || ((pixel_index >= 4586) && (pixel_index <= 4587)) || ((pixel_index >= 4589) && (pixel_index <= 4601)) || ((pixel_index >= 4613) && (pixel_index <= 4644)) || pixel_index == 4683 || ((pixel_index >= 4685) && (pixel_index <= 4697)) || ((pixel_index >= 4709) && (pixel_index <= 4742)) || ((pixel_index >= 4779) && (pixel_index <= 4793)) || ((pixel_index >= 4805) && (pixel_index <= 4838)) || ((pixel_index >= 4875) && (pixel_index <= 4889)) || ((pixel_index >= 4901) && (pixel_index <= 4934)) || ((pixel_index >= 4972) && (pixel_index <= 4985)) || ((pixel_index >= 4997) && (pixel_index <= 5029)) || ((pixel_index >= 5068) && (pixel_index <= 5081)) || ((pixel_index >= 5093) && (pixel_index <= 5125)) || ((pixel_index >= 5164) && (pixel_index <= 5177)) || ((pixel_index >= 5189) && (pixel_index <= 5221)) || ((pixel_index >= 5260) && (pixel_index <= 5273)) || ((pixel_index >= 5285) && (pixel_index <= 5316)) || ((pixel_index >= 5356) && (pixel_index <= 5369)) || ((pixel_index >= 5381) && (pixel_index <= 5412)) || ((pixel_index >= 5453) && (pixel_index <= 5465)) || ((pixel_index >= 5477) && (pixel_index <= 5508)) || ((pixel_index >= 5549) && (pixel_index <= 5561)) || ((pixel_index >= 5573) && (pixel_index <= 5604)) || ((pixel_index >= 5645) && (pixel_index <= 5649)) || ((pixel_index >= 5651) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5700)) || ((pixel_index >= 5741) && (pixel_index <= 5743)) || ((pixel_index >= 5747) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5796)) || ((pixel_index >= 5843) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5892)) || ((pixel_index >= 5937) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 5987)) || pixel_index == 6006 || ((pixel_index >= 6032) && (pixel_index <= 6041)) || ((pixel_index >= 6053) && (pixel_index <= 6083)) || pixel_index == 6102 || (pixel_index >= 6127) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 3) begin
            if (((pixel_index >= 5) && (pixel_index <= 56)) || ((pixel_index >= 68) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 152)) || ((pixel_index >= 164) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 248)) || ((pixel_index >= 261) && (pixel_index <= 262)) || ((pixel_index >= 264) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 345)) || ((pixel_index >= 363) && (pixel_index <= 377)) || ((pixel_index >= 389) && (pixel_index <= 441)) || ((pixel_index >= 460) && (pixel_index <= 473)) || ((pixel_index >= 485) && (pixel_index <= 534)) || ((pixel_index >= 557) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 628)) || ((pixel_index >= 653) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 722)) || ((pixel_index >= 750) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 817)) || ((pixel_index >= 846) && (pixel_index <= 857)) || ((pixel_index >= 869) && (pixel_index <= 912)) || ((pixel_index >= 942) && (pixel_index <= 953)) || ((pixel_index >= 965) && (pixel_index <= 1007)) || ((pixel_index >= 1039) && (pixel_index <= 1049)) || ((pixel_index >= 1061) && (pixel_index <= 1103)) || ((pixel_index >= 1135) && (pixel_index <= 1145)) || ((pixel_index >= 1157) && (pixel_index <= 1198)) || ((pixel_index >= 1232) && (pixel_index <= 1241)) || ((pixel_index >= 1253) && (pixel_index <= 1294)) || ((pixel_index >= 1328) && (pixel_index <= 1337)) || ((pixel_index >= 1349) && (pixel_index <= 1389)) || ((pixel_index >= 1424) && (pixel_index <= 1433)) || ((pixel_index >= 1445) && (pixel_index <= 1485)) || ((pixel_index >= 1521) && (pixel_index <= 1529)) || ((pixel_index >= 1541) && (pixel_index <= 1581)) || ((pixel_index >= 1617) && (pixel_index <= 1625)) || ((pixel_index >= 1637) && (pixel_index <= 1676)) || ((pixel_index >= 1713) && (pixel_index <= 1721)) || ((pixel_index >= 1733) && (pixel_index <= 1772)) || ((pixel_index >= 1810) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1869)) || ((pixel_index >= 1906) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 1965)) || ((pixel_index >= 2002) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2061)) || ((pixel_index >= 2098) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2158)) || ((pixel_index >= 2194) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2255)) || ((pixel_index >= 2291) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2352)) || ((pixel_index >= 2387) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2450)) || ((pixel_index >= 2483) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2546)) || ((pixel_index >= 2579) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2641)) || ((pixel_index >= 2675) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2737)) || ((pixel_index >= 2771) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2833)) || ((pixel_index >= 2867) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2930)) || ((pixel_index >= 2963) && (pixel_index <= 2969)) || ((pixel_index >= 2981) && (pixel_index <= 3027)) || ((pixel_index >= 3059) && (pixel_index <= 3065)) || ((pixel_index >= 3077) && (pixel_index <= 3124)) || ((pixel_index >= 3155) && (pixel_index <= 3161)) || ((pixel_index >= 3173) && (pixel_index <= 3207)) || ((pixel_index >= 3209) && (pixel_index <= 3210)) || ((pixel_index >= 3213) && (pixel_index <= 3220)) || ((pixel_index >= 3251) && (pixel_index <= 3257)) || ((pixel_index >= 3269) && (pixel_index <= 3302)) || ((pixel_index >= 3311) && (pixel_index <= 3317)) || ((pixel_index >= 3348) && (pixel_index <= 3353)) || ((pixel_index >= 3365) && (pixel_index <= 3396)) || ((pixel_index >= 3407) && (pixel_index <= 3414)) || ((pixel_index >= 3443) && (pixel_index <= 3449)) || ((pixel_index >= 3461) && (pixel_index <= 3491)) || ((pixel_index >= 3504) && (pixel_index <= 3510)) || ((pixel_index >= 3539) && (pixel_index <= 3545)) || ((pixel_index >= 3557) && (pixel_index <= 3586)) || ((pixel_index >= 3600) && (pixel_index <= 3605)) || ((pixel_index >= 3636) && (pixel_index <= 3641)) || ((pixel_index >= 3653) && (pixel_index <= 3682)) || ((pixel_index >= 3696) && (pixel_index <= 3702)) || ((pixel_index >= 3732) && (pixel_index <= 3737)) || ((pixel_index >= 3749) && (pixel_index <= 3778)) || ((pixel_index >= 3792) && (pixel_index <= 3798)) || ((pixel_index >= 3828) && (pixel_index <= 3833)) || ((pixel_index >= 3845) && (pixel_index <= 3874)) || ((pixel_index >= 3888) && (pixel_index <= 3894)) || ((pixel_index >= 3924) && (pixel_index <= 3929)) || ((pixel_index >= 3941) && (pixel_index <= 3970)) || ((pixel_index >= 3984) && (pixel_index <= 3991)) || pixel_index == 4015 || ((pixel_index >= 4020) && (pixel_index <= 4025)) || ((pixel_index >= 4037) && (pixel_index <= 4066)) || ((pixel_index >= 4080) && (pixel_index <= 4087)) || pixel_index == 4111 || pixel_index == 4114 || ((pixel_index >= 4116) && (pixel_index <= 4121)) || ((pixel_index >= 4133) && (pixel_index <= 4163)) || ((pixel_index >= 4177) && (pixel_index <= 4183)) || ((pixel_index >= 4207) && (pixel_index <= 4208)) || pixel_index == 4210 || ((pixel_index >= 4212) && (pixel_index <= 4217)) || ((pixel_index >= 4229) && (pixel_index <= 4259)) || ((pixel_index >= 4274) && (pixel_index <= 4279)) || ((pixel_index >= 4303) && (pixel_index <= 4304)) || ((pixel_index >= 4306) && (pixel_index <= 4313)) || ((pixel_index >= 4325) && (pixel_index <= 4356)) || ((pixel_index >= 4371) && (pixel_index <= 4375)) || ((pixel_index >= 4399) && (pixel_index <= 4409)) || ((pixel_index >= 4421) && (pixel_index <= 4452)) || ((pixel_index >= 4468) && (pixel_index <= 4470)) || ((pixel_index >= 4495) && (pixel_index <= 4505)) || ((pixel_index >= 4517) && (pixel_index <= 4549)) || ((pixel_index >= 4564) && (pixel_index <= 4566)) || ((pixel_index >= 4591) && (pixel_index <= 4601)) || ((pixel_index >= 4613) && (pixel_index <= 4647)) || pixel_index == 4661 || pixel_index == 4684 || ((pixel_index >= 4687) && (pixel_index <= 4697)) || ((pixel_index >= 4709) && (pixel_index <= 4743)) || ((pixel_index >= 4780) && (pixel_index <= 4781)) || ((pixel_index >= 4783) && (pixel_index <= 4793)) || ((pixel_index >= 4805) && (pixel_index <= 4839)) || ((pixel_index >= 4876) && (pixel_index <= 4889)) || ((pixel_index >= 4901) && (pixel_index <= 4935)) || ((pixel_index >= 4972) && (pixel_index <= 4985)) || ((pixel_index >= 4997) && (pixel_index <= 5030)) || ((pixel_index >= 5069) && (pixel_index <= 5081)) || ((pixel_index >= 5093) && (pixel_index <= 5126)) || ((pixel_index >= 5165) && (pixel_index <= 5177)) || ((pixel_index >= 5189) && (pixel_index <= 5222)) || ((pixel_index >= 5261) && (pixel_index <= 5273)) || ((pixel_index >= 5285) && (pixel_index <= 5317)) || ((pixel_index >= 5357) && (pixel_index <= 5369)) || ((pixel_index >= 5381) && (pixel_index <= 5413)) || ((pixel_index >= 5454) && (pixel_index <= 5465)) || ((pixel_index >= 5477) && (pixel_index <= 5509)) || ((pixel_index >= 5550) && (pixel_index <= 5561)) || ((pixel_index >= 5573) && (pixel_index <= 5605)) || ((pixel_index >= 5646) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5701)) || ((pixel_index >= 5742) && (pixel_index <= 5747)) || ((pixel_index >= 5749) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5797)) || ((pixel_index >= 5838) && (pixel_index <= 5841)) || ((pixel_index >= 5845) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5893)) || ((pixel_index >= 5935) && (pixel_index <= 5936)) || ((pixel_index >= 5941) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 5989)) || ((pixel_index >= 6036) && (pixel_index <= 6041)) || ((pixel_index >= 6053) && (pixel_index <= 6085)) || (pixel_index >= 6129) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 4) begin
            if (((pixel_index >= 5) && (pixel_index <= 57)) || ((pixel_index >= 69) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 153)) || ((pixel_index >= 166) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 250)) || ((pixel_index >= 266) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 346)) || ((pixel_index >= 364) && (pixel_index <= 377)) || ((pixel_index >= 389) && (pixel_index <= 439)) || ((pixel_index >= 461) && (pixel_index <= 473)) || ((pixel_index >= 485) && (pixel_index <= 533)) || ((pixel_index >= 558) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 627)) || ((pixel_index >= 654) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 722)) || ((pixel_index >= 751) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 817)) || ((pixel_index >= 847) && (pixel_index <= 857)) || ((pixel_index >= 869) && (pixel_index <= 912)) || ((pixel_index >= 944) && (pixel_index <= 953)) || ((pixel_index >= 965) && (pixel_index <= 1007)) || ((pixel_index >= 1040) && (pixel_index <= 1049)) || ((pixel_index >= 1061) && (pixel_index <= 1102)) || ((pixel_index >= 1136) && (pixel_index <= 1145)) || ((pixel_index >= 1157) && (pixel_index <= 1198)) || ((pixel_index >= 1233) && (pixel_index <= 1241)) || ((pixel_index >= 1253) && (pixel_index <= 1294)) || ((pixel_index >= 1329) && (pixel_index <= 1337)) || ((pixel_index >= 1349) && (pixel_index <= 1389)) || ((pixel_index >= 1425) && (pixel_index <= 1433)) || ((pixel_index >= 1445) && (pixel_index <= 1485)) || ((pixel_index >= 1522) && (pixel_index <= 1529)) || ((pixel_index >= 1541) && (pixel_index <= 1581)) || ((pixel_index >= 1618) && (pixel_index <= 1625)) || ((pixel_index >= 1637) && (pixel_index <= 1676)) || ((pixel_index >= 1714) && (pixel_index <= 1721)) || ((pixel_index >= 1733) && (pixel_index <= 1773)) || ((pixel_index >= 1810) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1869)) || ((pixel_index >= 1907) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 1965)) || ((pixel_index >= 2003) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2061)) || ((pixel_index >= 2099) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2158)) || ((pixel_index >= 2195) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2255)) || ((pixel_index >= 2292) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2352)) || ((pixel_index >= 2388) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2450)) || ((pixel_index >= 2484) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2546)) || ((pixel_index >= 2580) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2641)) || ((pixel_index >= 2676) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2736)) || ((pixel_index >= 2772) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2834)) || ((pixel_index >= 2868) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2930)) || ((pixel_index >= 2964) && (pixel_index <= 2969)) || ((pixel_index >= 2981) && (pixel_index <= 3027)) || ((pixel_index >= 3060) && (pixel_index <= 3065)) || ((pixel_index >= 3077) && (pixel_index <= 3113)) || ((pixel_index >= 3120) && (pixel_index <= 3124)) || ((pixel_index >= 3156) && (pixel_index <= 3161)) || ((pixel_index >= 3173) && (pixel_index <= 3206)) || ((pixel_index >= 3217) && (pixel_index <= 3220)) || ((pixel_index >= 3252) && (pixel_index <= 3257)) || ((pixel_index >= 3269) && (pixel_index <= 3301)) || ((pixel_index >= 3313) && (pixel_index <= 3317)) || ((pixel_index >= 3348) && (pixel_index <= 3353)) || ((pixel_index >= 3365) && (pixel_index <= 3396)) || ((pixel_index >= 3410) && (pixel_index <= 3414)) || ((pixel_index >= 3444) && (pixel_index <= 3449)) || ((pixel_index >= 3461) && (pixel_index <= 3492)) || ((pixel_index >= 3506) && (pixel_index <= 3510)) || ((pixel_index >= 3540) && (pixel_index <= 3545)) || ((pixel_index >= 3557) && (pixel_index <= 3588)) || ((pixel_index >= 3602) && (pixel_index <= 3606)) || ((pixel_index >= 3637) && (pixel_index <= 3641)) || ((pixel_index >= 3653) && (pixel_index <= 3683)) || ((pixel_index >= 3698) && (pixel_index <= 3702)) || ((pixel_index >= 3733) && (pixel_index <= 3737)) || ((pixel_index >= 3749) && (pixel_index <= 3779)) || ((pixel_index >= 3794) && (pixel_index <= 3798)) || ((pixel_index >= 3829) && (pixel_index <= 3833)) || ((pixel_index >= 3845) && (pixel_index <= 3876)) || ((pixel_index >= 3890) && (pixel_index <= 3895)) || ((pixel_index >= 3925) && (pixel_index <= 3929)) || ((pixel_index >= 3941) && (pixel_index <= 3972)) || ((pixel_index >= 3986) && (pixel_index <= 3991)) || ((pixel_index >= 4021) && (pixel_index <= 4025)) || ((pixel_index >= 4037) && (pixel_index <= 4068)) || ((pixel_index >= 4083) && (pixel_index <= 4087)) || ((pixel_index >= 4111) && (pixel_index <= 4112)) || ((pixel_index >= 4117) && (pixel_index <= 4121)) || ((pixel_index >= 4133) && (pixel_index <= 4164)) || ((pixel_index >= 4179) && (pixel_index <= 4183)) || pixel_index == 4208 || ((pixel_index >= 4213) && (pixel_index <= 4217)) || ((pixel_index >= 4229) && (pixel_index <= 4261)) || ((pixel_index >= 4276) && (pixel_index <= 4279)) || ((pixel_index >= 4304) && (pixel_index <= 4305)) || pixel_index == 4307 || ((pixel_index >= 4309) && (pixel_index <= 4313)) || ((pixel_index >= 4325) && (pixel_index <= 4358)) || ((pixel_index >= 4373) && (pixel_index <= 4375)) || ((pixel_index >= 4400) && (pixel_index <= 4401)) || ((pixel_index >= 4403) && (pixel_index <= 4409)) || ((pixel_index >= 4421) && (pixel_index <= 4455)) || pixel_index == 4470 || ((pixel_index >= 4496) && (pixel_index <= 4505)) || ((pixel_index >= 4517) && (pixel_index <= 4553)) || ((pixel_index >= 4592) && (pixel_index <= 4601)) || ((pixel_index >= 4613) && (pixel_index <= 4649)) || pixel_index == 4684 || ((pixel_index >= 4687) && (pixel_index <= 4697)) || ((pixel_index >= 4709) && (pixel_index <= 4744)) || ((pixel_index >= 4780) && (pixel_index <= 4781)) || ((pixel_index >= 4784) && (pixel_index <= 4793)) || ((pixel_index >= 4805) && (pixel_index <= 4840)) || ((pixel_index >= 4877) && (pixel_index <= 4878)) || ((pixel_index >= 4880) && (pixel_index <= 4889)) || ((pixel_index >= 4901) && (pixel_index <= 4935)) || ((pixel_index >= 4973) && (pixel_index <= 4974)) || ((pixel_index >= 4976) && (pixel_index <= 4985)) || ((pixel_index >= 4997) && (pixel_index <= 5031)) || ((pixel_index >= 5069) && (pixel_index <= 5081)) || ((pixel_index >= 5093) && (pixel_index <= 5127)) || ((pixel_index >= 5165) && (pixel_index <= 5177)) || ((pixel_index >= 5189) && (pixel_index <= 5223)) || ((pixel_index >= 5262) && (pixel_index <= 5273)) || ((pixel_index >= 5285) && (pixel_index <= 5319)) || ((pixel_index >= 5358) && (pixel_index <= 5369)) || ((pixel_index >= 5381) && (pixel_index <= 5415)) || ((pixel_index >= 5454) && (pixel_index <= 5465)) || ((pixel_index >= 5477) && (pixel_index <= 5511)) || ((pixel_index >= 5550) && (pixel_index <= 5561)) || ((pixel_index >= 5573) && (pixel_index <= 5607)) || ((pixel_index >= 5646) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5703)) || ((pixel_index >= 5743) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5798)) || ((pixel_index >= 5839) && (pixel_index <= 5843)) || ((pixel_index >= 5846) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5894)) || ((pixel_index >= 5935) && (pixel_index <= 5937)) || ((pixel_index >= 5942) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 5990)) || pixel_index == 6003 || ((pixel_index >= 6031) && (pixel_index <= 6032)) || ((pixel_index >= 6038) && (pixel_index <= 6041)) || ((pixel_index >= 6053) && (pixel_index <= 6086)) || ((pixel_index >= 6099) && (pixel_index <= 6100)) || (pixel_index >= 6132) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 5) begin
            if (((pixel_index >= 5) && (pixel_index <= 57)) || ((pixel_index >= 70) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 153)) || ((pixel_index >= 166) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 250)) || pixel_index == 263 || ((pixel_index >= 265) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 346)) || ((pixel_index >= 364) && (pixel_index <= 377)) || ((pixel_index >= 389) && (pixel_index <= 439)) || ((pixel_index >= 461) && (pixel_index <= 473)) || ((pixel_index >= 485) && (pixel_index <= 533)) || ((pixel_index >= 558) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 627)) || ((pixel_index >= 654) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 722)) || ((pixel_index >= 751) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 817)) || ((pixel_index >= 847) && (pixel_index <= 857)) || ((pixel_index >= 869) && (pixel_index <= 912)) || ((pixel_index >= 944) && (pixel_index <= 953)) || ((pixel_index >= 965) && (pixel_index <= 1007)) || ((pixel_index >= 1040) && (pixel_index <= 1049)) || ((pixel_index >= 1061) && (pixel_index <= 1102)) || ((pixel_index >= 1136) && (pixel_index <= 1145)) || ((pixel_index >= 1157) && (pixel_index <= 1198)) || ((pixel_index >= 1232) && (pixel_index <= 1241)) || ((pixel_index >= 1253) && (pixel_index <= 1294)) || ((pixel_index >= 1329) && (pixel_index <= 1337)) || ((pixel_index >= 1349) && (pixel_index <= 1389)) || ((pixel_index >= 1425) && (pixel_index <= 1433)) || ((pixel_index >= 1445) && (pixel_index <= 1485)) || ((pixel_index >= 1522) && (pixel_index <= 1529)) || ((pixel_index >= 1541) && (pixel_index <= 1580)) || ((pixel_index >= 1618) && (pixel_index <= 1625)) || ((pixel_index >= 1637) && (pixel_index <= 1676)) || ((pixel_index >= 1714) && (pixel_index <= 1721)) || ((pixel_index >= 1733) && (pixel_index <= 1772)) || ((pixel_index >= 1810) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1869)) || ((pixel_index >= 1907) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 1965)) || ((pixel_index >= 2003) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2061)) || ((pixel_index >= 2099) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2158)) || ((pixel_index >= 2195) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2255)) || ((pixel_index >= 2291) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2353)) || ((pixel_index >= 2388) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2449)) || ((pixel_index >= 2484) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2545)) || ((pixel_index >= 2580) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2640)) || ((pixel_index >= 2676) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2736)) || ((pixel_index >= 2772) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2833)) || ((pixel_index >= 2868) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2930)) || ((pixel_index >= 2964) && (pixel_index <= 2969)) || ((pixel_index >= 2981) && (pixel_index <= 3017)) || ((pixel_index >= 3019) && (pixel_index <= 3026)) || ((pixel_index >= 3060) && (pixel_index <= 3065)) || ((pixel_index >= 3077) && (pixel_index <= 3112)) || ((pixel_index >= 3121) && (pixel_index <= 3124)) || ((pixel_index >= 3156) && (pixel_index <= 3161)) || ((pixel_index >= 3173) && (pixel_index <= 3206)) || ((pixel_index >= 3218) && (pixel_index <= 3220)) || ((pixel_index >= 3252) && (pixel_index <= 3257)) || ((pixel_index >= 3269) && (pixel_index <= 3301)) || ((pixel_index >= 3314) && (pixel_index <= 3317)) || ((pixel_index >= 3348) && (pixel_index <= 3353)) || ((pixel_index >= 3365) && (pixel_index <= 3396)) || ((pixel_index >= 3410) && (pixel_index <= 3413)) || ((pixel_index >= 3444) && (pixel_index <= 3449)) || ((pixel_index >= 3461) && (pixel_index <= 3492)) || ((pixel_index >= 3506) && (pixel_index <= 3510)) || ((pixel_index >= 3540) && (pixel_index <= 3545)) || ((pixel_index >= 3557) && (pixel_index <= 3588)) || ((pixel_index >= 3603) && (pixel_index <= 3606)) || ((pixel_index >= 3637) && (pixel_index <= 3641)) || ((pixel_index >= 3653) && (pixel_index <= 3684)) || ((pixel_index >= 3698) && (pixel_index <= 3702)) || ((pixel_index >= 3733) && (pixel_index <= 3737)) || ((pixel_index >= 3749) && (pixel_index <= 3780)) || ((pixel_index >= 3794) && (pixel_index <= 3798)) || ((pixel_index >= 3829) && (pixel_index <= 3833)) || ((pixel_index >= 3845) && (pixel_index <= 3876)) || ((pixel_index >= 3890) && (pixel_index <= 3894)) || ((pixel_index >= 3925) && (pixel_index <= 3929)) || ((pixel_index >= 3941) && (pixel_index <= 3972)) || ((pixel_index >= 3987) && (pixel_index <= 3991)) || ((pixel_index >= 4021) && (pixel_index <= 4025)) || ((pixel_index >= 4037) && (pixel_index <= 4069)) || ((pixel_index >= 4084) && (pixel_index <= 4087)) || ((pixel_index >= 4111) && (pixel_index <= 4112)) || ((pixel_index >= 4117) && (pixel_index <= 4121)) || ((pixel_index >= 4133) && (pixel_index <= 4165)) || ((pixel_index >= 4180) && (pixel_index <= 4183)) || pixel_index == 4208 || ((pixel_index >= 4213) && (pixel_index <= 4217)) || ((pixel_index >= 4229) && (pixel_index <= 4262)) || ((pixel_index >= 4276) && (pixel_index <= 4279)) || pixel_index == 4304 || pixel_index == 4307 || ((pixel_index >= 4309) && (pixel_index <= 4313)) || ((pixel_index >= 4325) && (pixel_index <= 4359)) || ((pixel_index >= 4373) && (pixel_index <= 4375)) || ((pixel_index >= 4400) && (pixel_index <= 4401)) || ((pixel_index >= 4403) && (pixel_index <= 4409)) || ((pixel_index >= 4421) && (pixel_index <= 4456)) || pixel_index == 4470 || ((pixel_index >= 4496) && (pixel_index <= 4505)) || ((pixel_index >= 4517) && (pixel_index <= 4553)) || ((pixel_index >= 4592) && (pixel_index <= 4601)) || ((pixel_index >= 4613) && (pixel_index <= 4649)) || pixel_index == 4684 || ((pixel_index >= 4687) && (pixel_index <= 4697)) || ((pixel_index >= 4709) && (pixel_index <= 4744)) || ((pixel_index >= 4780) && (pixel_index <= 4781)) || ((pixel_index >= 4784) && (pixel_index <= 4793)) || ((pixel_index >= 4805) && (pixel_index <= 4840)) || ((pixel_index >= 4876) && (pixel_index <= 4878)) || ((pixel_index >= 4880) && (pixel_index <= 4889)) || ((pixel_index >= 4901) && (pixel_index <= 4936)) || ((pixel_index >= 4973) && (pixel_index <= 4974)) || ((pixel_index >= 4976) && (pixel_index <= 4985)) || ((pixel_index >= 4997) && (pixel_index <= 5032)) || ((pixel_index >= 5069) && (pixel_index <= 5070)) || ((pixel_index >= 5072) && (pixel_index <= 5081)) || ((pixel_index >= 5093) && (pixel_index <= 5128)) || ((pixel_index >= 5165) && (pixel_index <= 5177)) || ((pixel_index >= 5189) && (pixel_index <= 5223)) || ((pixel_index >= 5261) && (pixel_index <= 5273)) || ((pixel_index >= 5285) && (pixel_index <= 5319)) || ((pixel_index >= 5358) && (pixel_index <= 5369)) || ((pixel_index >= 5381) && (pixel_index <= 5415)) || ((pixel_index >= 5454) && (pixel_index <= 5465)) || ((pixel_index >= 5477) && (pixel_index <= 5511)) || ((pixel_index >= 5550) && (pixel_index <= 5561)) || ((pixel_index >= 5573) && (pixel_index <= 5606)) || ((pixel_index >= 5646) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5702)) || ((pixel_index >= 5743) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5798)) || ((pixel_index >= 5839) && (pixel_index <= 5843)) || ((pixel_index >= 5846) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5894)) || pixel_index == 5907 || ((pixel_index >= 5935) && (pixel_index <= 5937)) || ((pixel_index >= 5942) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 5990)) || pixel_index == 6003 || ((pixel_index >= 6031) && (pixel_index <= 6032)) || ((pixel_index >= 6037) && (pixel_index <= 6041)) || ((pixel_index >= 6053) && (pixel_index <= 6087)) || ((pixel_index >= 6098) && (pixel_index <= 6099)) || (pixel_index >= 6132) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
            done = 0;
        end
        else if (frame_count == 6) begin
            if (((pixel_index >= 5) && (pixel_index <= 57)) || ((pixel_index >= 70) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 153)) || ((pixel_index >= 166) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 250)) || ((pixel_index >= 263) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 346)) || ((pixel_index >= 363) && (pixel_index <= 377)) || ((pixel_index >= 389) && (pixel_index <= 440)) || ((pixel_index >= 461) && (pixel_index <= 473)) || ((pixel_index >= 485) && (pixel_index <= 533)) || ((pixel_index >= 557) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 627)) || ((pixel_index >= 654) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 722)) || ((pixel_index >= 751) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 817)) || ((pixel_index >= 847) && (pixel_index <= 857)) || ((pixel_index >= 869) && (pixel_index <= 912)) || ((pixel_index >= 943) && (pixel_index <= 953)) || ((pixel_index >= 965) && (pixel_index <= 1007)) || ((pixel_index >= 1040) && (pixel_index <= 1049)) || ((pixel_index >= 1061) && (pixel_index <= 1102)) || ((pixel_index >= 1136) && (pixel_index <= 1145)) || ((pixel_index >= 1157) && (pixel_index <= 1198)) || ((pixel_index >= 1232) && (pixel_index <= 1241)) || ((pixel_index >= 1253) && (pixel_index <= 1293)) || ((pixel_index >= 1329) && (pixel_index <= 1337)) || ((pixel_index >= 1349) && (pixel_index <= 1389)) || ((pixel_index >= 1425) && (pixel_index <= 1433)) || ((pixel_index >= 1445) && (pixel_index <= 1485)) || ((pixel_index >= 1521) && (pixel_index <= 1529)) || ((pixel_index >= 1541) && (pixel_index <= 1580)) || ((pixel_index >= 1618) && (pixel_index <= 1625)) || ((pixel_index >= 1637) && (pixel_index <= 1676)) || ((pixel_index >= 1714) && (pixel_index <= 1721)) || ((pixel_index >= 1733) && (pixel_index <= 1772)) || ((pixel_index >= 1810) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1868)) || ((pixel_index >= 1906) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 1965)) || ((pixel_index >= 2003) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2061)) || ((pixel_index >= 2099) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2158)) || ((pixel_index >= 2195) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2255)) || ((pixel_index >= 2291) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2352)) || ((pixel_index >= 2387) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2449)) || ((pixel_index >= 2484) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2545)) || ((pixel_index >= 2580) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2640)) || ((pixel_index >= 2676) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2736)) || ((pixel_index >= 2772) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2833)) || ((pixel_index >= 2868) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2929)) || ((pixel_index >= 2964) && (pixel_index <= 2969)) || ((pixel_index >= 2981) && (pixel_index <= 3017)) || pixel_index == 3019 || ((pixel_index >= 3021) && (pixel_index <= 3026)) || ((pixel_index >= 3060) && (pixel_index <= 3065)) || ((pixel_index >= 3077) && (pixel_index <= 3112)) || ((pixel_index >= 3121) && (pixel_index <= 3123)) || ((pixel_index >= 3156) && (pixel_index <= 3161)) || ((pixel_index >= 3173) && (pixel_index <= 3206)) || ((pixel_index >= 3217) && (pixel_index <= 3220)) || ((pixel_index >= 3252) && (pixel_index <= 3257)) || ((pixel_index >= 3269) && (pixel_index <= 3301)) || ((pixel_index >= 3314) && (pixel_index <= 3316)) || ((pixel_index >= 3348) && (pixel_index <= 3353)) || ((pixel_index >= 3365) && (pixel_index <= 3396)) || ((pixel_index >= 3410) && (pixel_index <= 3413)) || ((pixel_index >= 3444) && (pixel_index <= 3449)) || ((pixel_index >= 3461) && (pixel_index <= 3492)) || ((pixel_index >= 3506) && (pixel_index <= 3509)) || ((pixel_index >= 3540) && (pixel_index <= 3545)) || ((pixel_index >= 3557) && (pixel_index <= 3588)) || ((pixel_index >= 3602) && (pixel_index <= 3605)) || ((pixel_index >= 3636) && (pixel_index <= 3641)) || ((pixel_index >= 3653) && (pixel_index <= 3684)) || ((pixel_index >= 3698) && (pixel_index <= 3702)) || ((pixel_index >= 3732) && (pixel_index <= 3737)) || ((pixel_index >= 3749) && (pixel_index <= 3780)) || ((pixel_index >= 3794) && (pixel_index <= 3798)) || ((pixel_index >= 3829) && (pixel_index <= 3833)) || ((pixel_index >= 3845) && (pixel_index <= 3876)) || ((pixel_index >= 3890) && (pixel_index <= 3894)) || ((pixel_index >= 3925) && (pixel_index <= 3929)) || ((pixel_index >= 3941) && (pixel_index <= 3972)) || ((pixel_index >= 3987) && (pixel_index <= 3990)) || ((pixel_index >= 4021) && (pixel_index <= 4025)) || ((pixel_index >= 4037) && (pixel_index <= 4069)) || ((pixel_index >= 4083) && (pixel_index <= 4087)) || ((pixel_index >= 4117) && (pixel_index <= 4121)) || ((pixel_index >= 4133) && (pixel_index <= 4165)) || ((pixel_index >= 4180) && (pixel_index <= 4183)) || ((pixel_index >= 4207) && (pixel_index <= 4208)) || pixel_index == 4210 || ((pixel_index >= 4213) && (pixel_index <= 4217)) || ((pixel_index >= 4229) && (pixel_index <= 4262)) || ((pixel_index >= 4276) && (pixel_index <= 4279)) || pixel_index == 4304 || pixel_index == 4307 || ((pixel_index >= 4309) && (pixel_index <= 4313)) || ((pixel_index >= 4325) && (pixel_index <= 4359)) || ((pixel_index >= 4373) && (pixel_index <= 4375)) || ((pixel_index >= 4400) && (pixel_index <= 4401)) || pixel_index == 4403 || ((pixel_index >= 4405) && (pixel_index <= 4409)) || ((pixel_index >= 4421) && (pixel_index <= 4456)) || pixel_index == 4470 || ((pixel_index >= 4496) && (pixel_index <= 4497)) || ((pixel_index >= 4499) && (pixel_index <= 4505)) || ((pixel_index >= 4517) && (pixel_index <= 4553)) || ((pixel_index >= 4592) && (pixel_index <= 4601)) || ((pixel_index >= 4613) && (pixel_index <= 4649)) || pixel_index == 4684 || ((pixel_index >= 4687) && (pixel_index <= 4697)) || ((pixel_index >= 4709) && (pixel_index <= 4744)) || ((pixel_index >= 4780) && (pixel_index <= 4781)) || ((pixel_index >= 4784) && (pixel_index <= 4793)) || ((pixel_index >= 4805) && (pixel_index <= 4840)) || ((pixel_index >= 4876) && (pixel_index <= 4877)) || ((pixel_index >= 4880) && (pixel_index <= 4889)) || ((pixel_index >= 4901) && (pixel_index <= 4936)) || ((pixel_index >= 4973) && (pixel_index <= 4974)) || ((pixel_index >= 4976) && (pixel_index <= 4985)) || ((pixel_index >= 4997) && (pixel_index <= 5031)) || ((pixel_index >= 5069) && (pixel_index <= 5070)) || ((pixel_index >= 5072) && (pixel_index <= 5081)) || ((pixel_index >= 5093) && (pixel_index <= 5127)) || ((pixel_index >= 5165) && (pixel_index <= 5177)) || ((pixel_index >= 5189) && (pixel_index <= 5223)) || ((pixel_index >= 5261) && (pixel_index <= 5273)) || ((pixel_index >= 5285) && (pixel_index <= 5319)) || ((pixel_index >= 5358) && (pixel_index <= 5369)) || ((pixel_index >= 5381) && (pixel_index <= 5415)) || ((pixel_index >= 5454) && (pixel_index <= 5465)) || ((pixel_index >= 5477) && (pixel_index <= 5510)) || ((pixel_index >= 5550) && (pixel_index <= 5561)) || ((pixel_index >= 5573) && (pixel_index <= 5606)) || ((pixel_index >= 5646) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5702)) || ((pixel_index >= 5743) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5798)) || pixel_index == 5811 || ((pixel_index >= 5839) && (pixel_index <= 5843)) || ((pixel_index >= 5846) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5894)) || ((pixel_index >= 5906) && (pixel_index <= 5907)) || ((pixel_index >= 5935) && (pixel_index <= 5937)) || ((pixel_index >= 5942) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 5990)) || ((pixel_index >= 6002) && (pixel_index <= 6003)) || pixel_index == 6031 || ((pixel_index >= 6037) && (pixel_index <= 6041)) || ((pixel_index >= 6053) && (pixel_index <= 6086)) || ((pixel_index >= 6097) && (pixel_index <= 6099)) || (pixel_index >= 6131) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 7) begin
            if (((pixel_index >= 5) && (pixel_index <= 57)) || ((pixel_index >= 69) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 153)) || ((pixel_index >= 166) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 249)) || ((pixel_index >= 262) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 346)) || ((pixel_index >= 363) && (pixel_index <= 377)) || ((pixel_index >= 389) && (pixel_index <= 439)) || ((pixel_index >= 460) && (pixel_index <= 473)) || ((pixel_index >= 485) && (pixel_index <= 533)) || ((pixel_index >= 557) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 627)) || ((pixel_index >= 654) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 722)) || ((pixel_index >= 750) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 816)) || ((pixel_index >= 847) && (pixel_index <= 857)) || ((pixel_index >= 869) && (pixel_index <= 911)) || ((pixel_index >= 943) && (pixel_index <= 953)) || ((pixel_index >= 965) && (pixel_index <= 1007)) || ((pixel_index >= 1039) && (pixel_index <= 1049)) || ((pixel_index >= 1061) && (pixel_index <= 1102)) || ((pixel_index >= 1135) && (pixel_index <= 1145)) || ((pixel_index >= 1157) && (pixel_index <= 1197)) || ((pixel_index >= 1232) && (pixel_index <= 1241)) || ((pixel_index >= 1253) && (pixel_index <= 1293)) || ((pixel_index >= 1328) && (pixel_index <= 1337)) || ((pixel_index >= 1349) && (pixel_index <= 1389)) || ((pixel_index >= 1425) && (pixel_index <= 1433)) || ((pixel_index >= 1445) && (pixel_index <= 1484)) || ((pixel_index >= 1521) && (pixel_index <= 1529)) || ((pixel_index >= 1541) && (pixel_index <= 1580)) || ((pixel_index >= 1617) && (pixel_index <= 1625)) || ((pixel_index >= 1637) && (pixel_index <= 1676)) || ((pixel_index >= 1714) && (pixel_index <= 1721)) || ((pixel_index >= 1733) && (pixel_index <= 1772)) || ((pixel_index >= 1810) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1868)) || ((pixel_index >= 1906) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 1964)) || ((pixel_index >= 2002) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2061)) || ((pixel_index >= 2099) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2157)) || ((pixel_index >= 2195) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2254)) || ((pixel_index >= 2291) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2352)) || ((pixel_index >= 2387) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2449)) || ((pixel_index >= 2483) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2545)) || ((pixel_index >= 2579) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2640)) || ((pixel_index >= 2675) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2735)) || ((pixel_index >= 2772) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2833)) || ((pixel_index >= 2868) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2929)) || ((pixel_index >= 2964) && (pixel_index <= 2969)) || ((pixel_index >= 2981) && (pixel_index <= 3025)) || ((pixel_index >= 3060) && (pixel_index <= 3065)) || ((pixel_index >= 3077) && (pixel_index <= 3112)) || ((pixel_index >= 3120) && (pixel_index <= 3123)) || ((pixel_index >= 3156) && (pixel_index <= 3161)) || ((pixel_index >= 3173) && (pixel_index <= 3206)) || ((pixel_index >= 3217) && (pixel_index <= 3219)) || ((pixel_index >= 3252) && (pixel_index <= 3257)) || ((pixel_index >= 3269) && (pixel_index <= 3301)) || ((pixel_index >= 3313) && (pixel_index <= 3316)) || ((pixel_index >= 3348) && (pixel_index <= 3353)) || ((pixel_index >= 3365) && (pixel_index <= 3396)) || ((pixel_index >= 3410) && (pixel_index <= 3413)) || ((pixel_index >= 3444) && (pixel_index <= 3449)) || ((pixel_index >= 3461) && (pixel_index <= 3492)) || ((pixel_index >= 3506) && (pixel_index <= 3509)) || ((pixel_index >= 3540) && (pixel_index <= 3545)) || ((pixel_index >= 3557) && (pixel_index <= 3587)) || ((pixel_index >= 3602) && (pixel_index <= 3605)) || ((pixel_index >= 3636) && (pixel_index <= 3641)) || ((pixel_index >= 3653) && (pixel_index <= 3683)) || ((pixel_index >= 3698) && (pixel_index <= 3701)) || ((pixel_index >= 3732) && (pixel_index <= 3737)) || ((pixel_index >= 3749) && (pixel_index <= 3779)) || ((pixel_index >= 3794) && (pixel_index <= 3798)) || ((pixel_index >= 3828) && (pixel_index <= 3833)) || ((pixel_index >= 3845) && (pixel_index <= 3876)) || ((pixel_index >= 3890) && (pixel_index <= 3894)) || ((pixel_index >= 3924) && (pixel_index <= 3929)) || ((pixel_index >= 3941) && (pixel_index <= 3972)) || ((pixel_index >= 3986) && (pixel_index <= 3990)) || pixel_index == 4015 || ((pixel_index >= 4020) && (pixel_index <= 4025)) || ((pixel_index >= 4037) && (pixel_index <= 4068)) || ((pixel_index >= 4083) && (pixel_index <= 4086)) || pixel_index == 4111 || ((pixel_index >= 4116) && (pixel_index <= 4121)) || ((pixel_index >= 4133) && (pixel_index <= 4165)) || ((pixel_index >= 4179) && (pixel_index <= 4183)) || ((pixel_index >= 4207) && (pixel_index <= 4208)) || pixel_index == 4210 || ((pixel_index >= 4213) && (pixel_index <= 4217)) || ((pixel_index >= 4229) && (pixel_index <= 4261)) || ((pixel_index >= 4276) && (pixel_index <= 4279)) || pixel_index == 4304 || ((pixel_index >= 4306) && (pixel_index <= 4307)) || ((pixel_index >= 4309) && (pixel_index <= 4313)) || ((pixel_index >= 4325) && (pixel_index <= 4358)) || ((pixel_index >= 4373) && (pixel_index <= 4375)) || ((pixel_index >= 4400) && (pixel_index <= 4403)) || ((pixel_index >= 4405) && (pixel_index <= 4409)) || ((pixel_index >= 4421) && (pixel_index <= 4455)) || pixel_index == 4470 || ((pixel_index >= 4496) && (pixel_index <= 4497)) || ((pixel_index >= 4499) && (pixel_index <= 4505)) || ((pixel_index >= 4517) && (pixel_index <= 4553)) || ((pixel_index >= 4591) && (pixel_index <= 4601)) || ((pixel_index >= 4613) && (pixel_index <= 4648)) || ((pixel_index >= 4687) && (pixel_index <= 4697)) || ((pixel_index >= 4709) && (pixel_index <= 4744)) || pixel_index == 4780 || ((pixel_index >= 4783) && (pixel_index <= 4793)) || ((pixel_index >= 4805) && (pixel_index <= 4839)) || ((pixel_index >= 4876) && (pixel_index <= 4877)) || ((pixel_index >= 4879) && (pixel_index <= 4889)) || ((pixel_index >= 4901) && (pixel_index <= 4935)) || ((pixel_index >= 4973) && (pixel_index <= 4974)) || ((pixel_index >= 4976) && (pixel_index <= 4985)) || ((pixel_index >= 4997) && (pixel_index <= 5031)) || ((pixel_index >= 5069) && (pixel_index <= 5070)) || ((pixel_index >= 5072) && (pixel_index <= 5081)) || ((pixel_index >= 5093) && (pixel_index <= 5127)) || ((pixel_index >= 5165) && (pixel_index <= 5177)) || ((pixel_index >= 5189) && (pixel_index <= 5223)) || ((pixel_index >= 5261) && (pixel_index <= 5273)) || ((pixel_index >= 5285) && (pixel_index <= 5318)) || ((pixel_index >= 5358) && (pixel_index <= 5369)) || ((pixel_index >= 5381) && (pixel_index <= 5414)) || ((pixel_index >= 5454) && (pixel_index <= 5465)) || ((pixel_index >= 5477) && (pixel_index <= 5510)) || ((pixel_index >= 5550) && (pixel_index <= 5561)) || ((pixel_index >= 5573) && (pixel_index <= 5606)) || ((pixel_index >= 5646) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5702)) || pixel_index == 5715 || ((pixel_index >= 5743) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5798)) || pixel_index == 5811 || ((pixel_index >= 5839) && (pixel_index <= 5843)) || ((pixel_index >= 5846) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5894)) || ((pixel_index >= 5906) && (pixel_index <= 5907)) || ((pixel_index >= 5935) && (pixel_index <= 5937)) || ((pixel_index >= 5942) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 5990)) || ((pixel_index >= 6001) && (pixel_index <= 6003)) || ((pixel_index >= 6031) && (pixel_index <= 6032)) || ((pixel_index >= 6037) && (pixel_index <= 6041)) || ((pixel_index >= 6053) && (pixel_index <= 6086)) || ((pixel_index >= 6097) && (pixel_index <= 6099)) || (pixel_index >= 6131) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 8) begin
            if (((pixel_index >= 5) && (pixel_index <= 55)) || ((pixel_index >= 68) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 151)) || ((pixel_index >= 165) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 248)) || ((pixel_index >= 264) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 345)) || ((pixel_index >= 362) && (pixel_index <= 377)) || ((pixel_index >= 389) && (pixel_index <= 440)) || ((pixel_index >= 459) && (pixel_index <= 473)) || ((pixel_index >= 485) && (pixel_index <= 533)) || ((pixel_index >= 556) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 627)) || ((pixel_index >= 653) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 721)) || ((pixel_index >= 749) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 816)) || ((pixel_index >= 846) && (pixel_index <= 857)) || ((pixel_index >= 869) && (pixel_index <= 911)) || ((pixel_index >= 942) && (pixel_index <= 953)) || ((pixel_index >= 965) && (pixel_index <= 1006)) || ((pixel_index >= 1039) && (pixel_index <= 1049)) || ((pixel_index >= 1061) && (pixel_index <= 1102)) || ((pixel_index >= 1135) && (pixel_index <= 1145)) || ((pixel_index >= 1157) && (pixel_index <= 1197)) || ((pixel_index >= 1231) && (pixel_index <= 1241)) || ((pixel_index >= 1253) && (pixel_index <= 1293)) || ((pixel_index >= 1328) && (pixel_index <= 1337)) || ((pixel_index >= 1349) && (pixel_index <= 1388)) || ((pixel_index >= 1424) && (pixel_index <= 1433)) || ((pixel_index >= 1445) && (pixel_index <= 1484)) || ((pixel_index >= 1521) && (pixel_index <= 1529)) || ((pixel_index >= 1541) && (pixel_index <= 1580)) || ((pixel_index >= 1617) && (pixel_index <= 1625)) || ((pixel_index >= 1637) && (pixel_index <= 1675)) || ((pixel_index >= 1713) && (pixel_index <= 1721)) || ((pixel_index >= 1733) && (pixel_index <= 1771)) || ((pixel_index >= 1809) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1867)) || ((pixel_index >= 1906) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 1964)) || ((pixel_index >= 2002) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2060)) || ((pixel_index >= 2098) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2156)) || ((pixel_index >= 2194) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2253)) || ((pixel_index >= 2291) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2350)) || ((pixel_index >= 2387) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2448)) || ((pixel_index >= 2483) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2545)) || ((pixel_index >= 2579) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2640)) || ((pixel_index >= 2675) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2736)) || ((pixel_index >= 2771) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2832)) || ((pixel_index >= 2867) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2929)) || ((pixel_index >= 2963) && (pixel_index <= 2969)) || ((pixel_index >= 2981) && (pixel_index <= 3025)) || ((pixel_index >= 3059) && (pixel_index <= 3065)) || ((pixel_index >= 3077) && (pixel_index <= 3122)) || ((pixel_index >= 3155) && (pixel_index <= 3161)) || ((pixel_index >= 3173) && (pixel_index <= 3207)) || ((pixel_index >= 3215) && (pixel_index <= 3219)) || ((pixel_index >= 3252) && (pixel_index <= 3257)) || ((pixel_index >= 3269) && (pixel_index <= 3301)) || ((pixel_index >= 3312) && (pixel_index <= 3316)) || ((pixel_index >= 3348) && (pixel_index <= 3353)) || ((pixel_index >= 3365) && (pixel_index <= 3396)) || ((pixel_index >= 3408) && (pixel_index <= 3412)) || ((pixel_index >= 3444) && (pixel_index <= 3449)) || ((pixel_index >= 3461) && (pixel_index <= 3491)) || ((pixel_index >= 3505) && (pixel_index <= 3509)) || ((pixel_index >= 3540) && (pixel_index <= 3545)) || ((pixel_index >= 3557) && (pixel_index <= 3587)) || ((pixel_index >= 3601) && (pixel_index <= 3605)) || ((pixel_index >= 3636) && (pixel_index <= 3641)) || ((pixel_index >= 3653) && (pixel_index <= 3682)) || ((pixel_index >= 3697) && (pixel_index <= 3701)) || ((pixel_index >= 3732) && (pixel_index <= 3737)) || ((pixel_index >= 3749) && (pixel_index <= 3778)) || ((pixel_index >= 3793) && (pixel_index <= 3797)) || ((pixel_index >= 3828) && (pixel_index <= 3833)) || ((pixel_index >= 3845) && (pixel_index <= 3874)) || ((pixel_index >= 3889) && (pixel_index <= 3894)) || ((pixel_index >= 3924) && (pixel_index <= 3929)) || ((pixel_index >= 3941) && (pixel_index <= 3971)) || ((pixel_index >= 3985) && (pixel_index <= 3990)) || pixel_index == 4015 || ((pixel_index >= 4020) && (pixel_index <= 4025)) || ((pixel_index >= 4037) && (pixel_index <= 4067)) || ((pixel_index >= 4082) && (pixel_index <= 4086)) || pixel_index == 4111 || ((pixel_index >= 4116) && (pixel_index <= 4121)) || ((pixel_index >= 4133) && (pixel_index <= 4163)) || ((pixel_index >= 4178) && (pixel_index <= 4182)) || ((pixel_index >= 4207) && (pixel_index <= 4208)) || pixel_index == 4210 || ((pixel_index >= 4212) && (pixel_index <= 4217)) || ((pixel_index >= 4229) && (pixel_index <= 4260)) || ((pixel_index >= 4275) && (pixel_index <= 4278)) || ((pixel_index >= 4303) && (pixel_index <= 4304)) || ((pixel_index >= 4306) && (pixel_index <= 4313)) || ((pixel_index >= 4325) && (pixel_index <= 4356)) || ((pixel_index >= 4372) && (pixel_index <= 4375)) || ((pixel_index >= 4399) && (pixel_index <= 4409)) || ((pixel_index >= 4421) && (pixel_index <= 4453)) || ((pixel_index >= 4468) && (pixel_index <= 4470)) || ((pixel_index >= 4495) && (pixel_index <= 4505)) || ((pixel_index >= 4517) && (pixel_index <= 4550)) || ((pixel_index >= 4591) && (pixel_index <= 4601)) || ((pixel_index >= 4613) && (pixel_index <= 4648)) || ((pixel_index >= 4687) && (pixel_index <= 4697)) || ((pixel_index >= 4709) && (pixel_index <= 4743)) || ((pixel_index >= 4780) && (pixel_index <= 4781)) || ((pixel_index >= 4783) && (pixel_index <= 4793)) || ((pixel_index >= 4805) && (pixel_index <= 4839)) || pixel_index == 4877 || ((pixel_index >= 4879) && (pixel_index <= 4889)) || ((pixel_index >= 4901) && (pixel_index <= 4935)) || ((pixel_index >= 4973) && (pixel_index <= 4985)) || ((pixel_index >= 4997) && (pixel_index <= 5030)) || ((pixel_index >= 5069) && (pixel_index <= 5081)) || ((pixel_index >= 5093) && (pixel_index <= 5126)) || ((pixel_index >= 5165) && (pixel_index <= 5177)) || ((pixel_index >= 5189) && (pixel_index <= 5222)) || ((pixel_index >= 5262) && (pixel_index <= 5273)) || ((pixel_index >= 5285) && (pixel_index <= 5318)) || ((pixel_index >= 5358) && (pixel_index <= 5369)) || ((pixel_index >= 5381) && (pixel_index <= 5414)) || ((pixel_index >= 5454) && (pixel_index <= 5465)) || ((pixel_index >= 5477) && (pixel_index <= 5510)) || ((pixel_index >= 5550) && (pixel_index <= 5561)) || ((pixel_index >= 5573) && (pixel_index <= 5606)) || ((pixel_index >= 5646) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5702)) || pixel_index == 5715 || ((pixel_index >= 5743) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5798)) || pixel_index == 5811 || ((pixel_index >= 5839) && (pixel_index <= 5844)) || ((pixel_index >= 5847) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5893)) || ((pixel_index >= 5906) && (pixel_index <= 5907)) || ((pixel_index >= 5935) && (pixel_index <= 5938)) || ((pixel_index >= 5943) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 5989)) || ((pixel_index >= 6001) && (pixel_index <= 6003)) || pixel_index == 6032 || ((pixel_index >= 6038) && (pixel_index <= 6041)) || ((pixel_index >= 6053) && (pixel_index <= 6085)) || ((pixel_index >= 6097) && (pixel_index <= 6099)) || (pixel_index >= 6132) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 9) begin
            if (((pixel_index >= 5) && (pixel_index <= 52)) || ((pixel_index >= 65) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 148)) || ((pixel_index >= 161) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 244)) || ((pixel_index >= 263) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 341)) || ((pixel_index >= 361) && (pixel_index <= 377)) || ((pixel_index >= 389) && (pixel_index <= 438)) || ((pixel_index >= 458) && (pixel_index <= 473)) || ((pixel_index >= 485) && (pixel_index <= 532)) || ((pixel_index >= 554) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 626)) || ((pixel_index >= 651) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 720)) || ((pixel_index >= 748) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 815)) || ((pixel_index >= 844) && (pixel_index <= 857)) || ((pixel_index >= 869) && (pixel_index <= 910)) || ((pixel_index >= 940) && (pixel_index <= 953)) || ((pixel_index >= 965) && (pixel_index <= 1005)) || ((pixel_index >= 1037) && (pixel_index <= 1049)) || ((pixel_index >= 1061) && (pixel_index <= 1100)) || ((pixel_index >= 1133) && (pixel_index <= 1145)) || ((pixel_index >= 1157) && (pixel_index <= 1196)) || ((pixel_index >= 1230) && (pixel_index <= 1241)) || ((pixel_index >= 1253) && (pixel_index <= 1291)) || ((pixel_index >= 1326) && (pixel_index <= 1337)) || ((pixel_index >= 1349) && (pixel_index <= 1387)) || ((pixel_index >= 1423) && (pixel_index <= 1433)) || ((pixel_index >= 1445) && (pixel_index <= 1482)) || ((pixel_index >= 1519) && (pixel_index <= 1529)) || ((pixel_index >= 1541) && (pixel_index <= 1578)) || ((pixel_index >= 1615) && (pixel_index <= 1625)) || ((pixel_index >= 1637) && (pixel_index <= 1674)) || ((pixel_index >= 1712) && (pixel_index <= 1721)) || ((pixel_index >= 1733) && (pixel_index <= 1770)) || ((pixel_index >= 1808) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1865)) || ((pixel_index >= 1904) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 1962)) || ((pixel_index >= 2001) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2058)) || ((pixel_index >= 2097) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2154)) || ((pixel_index >= 2193) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2250)) || ((pixel_index >= 2289) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2347)) || ((pixel_index >= 2385) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2444)) || ((pixel_index >= 2482) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2542)) || ((pixel_index >= 2578) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2639)) || ((pixel_index >= 2674) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2735)) || ((pixel_index >= 2770) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2831)) || ((pixel_index >= 2866) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2926)) || ((pixel_index >= 2962) && (pixel_index <= 2969)) || ((pixel_index >= 2981) && (pixel_index <= 3024)) || ((pixel_index >= 3058) && (pixel_index <= 3065)) || ((pixel_index >= 3077) && (pixel_index <= 3120)) || ((pixel_index >= 3154) && (pixel_index <= 3161)) || ((pixel_index >= 3173) && (pixel_index <= 3210)) || ((pixel_index >= 3212) && (pixel_index <= 3217)) || ((pixel_index >= 3250) && (pixel_index <= 3257)) || ((pixel_index >= 3269) && (pixel_index <= 3302)) || ((pixel_index >= 3310) && (pixel_index <= 3314)) || ((pixel_index >= 3347) && (pixel_index <= 3353)) || ((pixel_index >= 3365) && (pixel_index <= 3395)) || ((pixel_index >= 3407) && (pixel_index <= 3411)) || ((pixel_index >= 3443) && (pixel_index <= 3449)) || ((pixel_index >= 3461) && (pixel_index <= 3490)) || ((pixel_index >= 3503) && (pixel_index <= 3508)) || ((pixel_index >= 3539) && (pixel_index <= 3545)) || ((pixel_index >= 3557) && (pixel_index <= 3586)) || ((pixel_index >= 3599) && (pixel_index <= 3604)) || ((pixel_index >= 3635) && (pixel_index <= 3641)) || ((pixel_index >= 3653) && (pixel_index <= 3681)) || ((pixel_index >= 3696) && (pixel_index <= 3700)) || ((pixel_index >= 3731) && (pixel_index <= 3737)) || ((pixel_index >= 3749) && (pixel_index <= 3777)) || ((pixel_index >= 3792) && (pixel_index <= 3796)) || ((pixel_index >= 3827) && (pixel_index <= 3833)) || ((pixel_index >= 3845) && (pixel_index <= 3873)) || ((pixel_index >= 3887) && (pixel_index <= 3893)) || ((pixel_index >= 3923) && (pixel_index <= 3929)) || ((pixel_index >= 3941) && (pixel_index <= 3969)) || ((pixel_index >= 3983) && (pixel_index <= 3989)) || pixel_index == 4014 || ((pixel_index >= 4019) && (pixel_index <= 4025)) || ((pixel_index >= 4037) && (pixel_index <= 4065)) || ((pixel_index >= 4080) && (pixel_index <= 4085)) || pixel_index == 4110 || ((pixel_index >= 4115) && (pixel_index <= 4121)) || ((pixel_index >= 4133) && (pixel_index <= 4162)) || ((pixel_index >= 4177) && (pixel_index <= 4181)) || ((pixel_index >= 4206) && (pixel_index <= 4207)) || pixel_index == 4209 || ((pixel_index >= 4212) && (pixel_index <= 4217)) || ((pixel_index >= 4229) && (pixel_index <= 4258)) || ((pixel_index >= 4273) && (pixel_index <= 4277)) || ((pixel_index >= 4302) && (pixel_index <= 4303)) || ((pixel_index >= 4305) && (pixel_index <= 4306)) || ((pixel_index >= 4308) && (pixel_index <= 4313)) || ((pixel_index >= 4325) && (pixel_index <= 4354)) || ((pixel_index >= 4370) && (pixel_index <= 4374)) || ((pixel_index >= 4399) && (pixel_index <= 4409)) || ((pixel_index >= 4421) && (pixel_index <= 4451)) || ((pixel_index >= 4467) && (pixel_index <= 4469)) || ((pixel_index >= 4494) && (pixel_index <= 4505)) || ((pixel_index >= 4517) && (pixel_index <= 4548)) || ((pixel_index >= 4563) && (pixel_index <= 4564)) || ((pixel_index >= 4590) && (pixel_index <= 4601)) || ((pixel_index >= 4613) && (pixel_index <= 4645)) || ((pixel_index >= 4686) && (pixel_index <= 4697)) || ((pixel_index >= 4709) && (pixel_index <= 4743)) || pixel_index == 4780 || ((pixel_index >= 4783) && (pixel_index <= 4793)) || ((pixel_index >= 4805) && (pixel_index <= 4838)) || ((pixel_index >= 4876) && (pixel_index <= 4877)) || ((pixel_index >= 4879) && (pixel_index <= 4889)) || ((pixel_index >= 4901) && (pixel_index <= 4934)) || ((pixel_index >= 4972) && (pixel_index <= 4973)) || ((pixel_index >= 4975) && (pixel_index <= 4985)) || ((pixel_index >= 4997) && (pixel_index <= 5029)) || ((pixel_index >= 5068) && (pixel_index <= 5081)) || ((pixel_index >= 5093) && (pixel_index <= 5125)) || ((pixel_index >= 5165) && (pixel_index <= 5177)) || ((pixel_index >= 5189) && (pixel_index <= 5221)) || ((pixel_index >= 5261) && (pixel_index <= 5273)) || ((pixel_index >= 5285) && (pixel_index <= 5317)) || ((pixel_index >= 5357) && (pixel_index <= 5369)) || ((pixel_index >= 5381) && (pixel_index <= 5413)) || ((pixel_index >= 5454) && (pixel_index <= 5465)) || ((pixel_index >= 5477) && (pixel_index <= 5509)) || ((pixel_index >= 5550) && (pixel_index <= 5561)) || ((pixel_index >= 5573) && (pixel_index <= 5605)) || ((pixel_index >= 5646) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5701)) || ((pixel_index >= 5742) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5797)) || pixel_index == 5810 || ((pixel_index >= 5839) && (pixel_index <= 5843)) || ((pixel_index >= 5847) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5892)) || pixel_index == 5906 || ((pixel_index >= 5935) && (pixel_index <= 5938)) || ((pixel_index >= 5942) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 5988)) || ((pixel_index >= 6001) && (pixel_index <= 6002)) || pixel_index == 6032 || ((pixel_index >= 6038) && (pixel_index <= 6041)) || ((pixel_index >= 6053) && (pixel_index <= 6084)) || ((pixel_index >= 6097) && (pixel_index <= 6098)) || (pixel_index >= 6132) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 10) begin
            if (((pixel_index >= 5) && (pixel_index <= 47)) || ((pixel_index >= 61) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 143)) || ((pixel_index >= 158) && (pixel_index <= 160)) || ((pixel_index >= 163) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 240)) || ((pixel_index >= 262) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 336)) || ((pixel_index >= 359) && (pixel_index <= 377)) || ((pixel_index >= 389) && (pixel_index <= 433)) || ((pixel_index >= 456) && (pixel_index <= 473)) || ((pixel_index >= 485) && (pixel_index <= 530)) || ((pixel_index >= 553) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 625)) || ((pixel_index >= 649) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 719)) || ((pixel_index >= 746) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 814)) || ((pixel_index >= 842) && (pixel_index <= 857)) || ((pixel_index >= 869) && (pixel_index <= 909)) || ((pixel_index >= 938) && (pixel_index <= 953)) || ((pixel_index >= 965) && (pixel_index <= 1004)) || ((pixel_index >= 1035) && (pixel_index <= 1049)) || ((pixel_index >= 1061) && (pixel_index <= 1099)) || ((pixel_index >= 1131) && (pixel_index <= 1145)) || ((pixel_index >= 1157) && (pixel_index <= 1194)) || ((pixel_index >= 1227) && (pixel_index <= 1241)) || ((pixel_index >= 1253) && (pixel_index <= 1290)) || ((pixel_index >= 1324) && (pixel_index <= 1337)) || ((pixel_index >= 1349) && (pixel_index <= 1385)) || ((pixel_index >= 1420) && (pixel_index <= 1433)) || ((pixel_index >= 1445) && (pixel_index <= 1481)) || ((pixel_index >= 1517) && (pixel_index <= 1529)) || ((pixel_index >= 1541) && (pixel_index <= 1577)) || ((pixel_index >= 1613) && (pixel_index <= 1625)) || ((pixel_index >= 1637) && (pixel_index <= 1673)) || ((pixel_index >= 1709) && (pixel_index <= 1721)) || ((pixel_index >= 1733) && (pixel_index <= 1768)) || ((pixel_index >= 1806) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1864)) || ((pixel_index >= 1902) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 1960)) || ((pixel_index >= 1998) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2056)) || ((pixel_index >= 2094) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2152)) || ((pixel_index >= 2191) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2249)) || ((pixel_index >= 2287) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2345)) || ((pixel_index >= 2383) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2442)) || ((pixel_index >= 2479) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2539)) || ((pixel_index >= 2575) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2638)) || ((pixel_index >= 2671) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2735)) || ((pixel_index >= 2767) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2831)) || ((pixel_index >= 2863) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2926)) || ((pixel_index >= 2960) && (pixel_index <= 2969)) || ((pixel_index >= 2981) && (pixel_index <= 3022)) || ((pixel_index >= 3056) && (pixel_index <= 3065)) || ((pixel_index >= 3077) && (pixel_index <= 3119)) || ((pixel_index >= 3152) && (pixel_index <= 3161)) || ((pixel_index >= 3173) && (pixel_index <= 3216)) || ((pixel_index >= 3248) && (pixel_index <= 3257)) || ((pixel_index >= 3269) && (pixel_index <= 3313)) || ((pixel_index >= 3344) && (pixel_index <= 3353)) || ((pixel_index >= 3365) && (pixel_index <= 3396)) || ((pixel_index >= 3404) && (pixel_index <= 3410)) || ((pixel_index >= 3440) && (pixel_index <= 3449)) || ((pixel_index >= 3461) && (pixel_index <= 3490)) || ((pixel_index >= 3501) && (pixel_index <= 3506)) || pixel_index == 3512 || ((pixel_index >= 3536) && (pixel_index <= 3545)) || ((pixel_index >= 3557) && (pixel_index <= 3585)) || ((pixel_index >= 3597) && (pixel_index <= 3602)) || ((pixel_index >= 3608) && (pixel_index <= 3609)) || ((pixel_index >= 3632) && (pixel_index <= 3641)) || ((pixel_index >= 3653) && (pixel_index <= 3680)) || ((pixel_index >= 3693) && (pixel_index <= 3698)) || ((pixel_index >= 3704) && (pixel_index <= 3705)) || ((pixel_index >= 3728) && (pixel_index <= 3737)) || ((pixel_index >= 3749) && (pixel_index <= 3776)) || ((pixel_index >= 3790) && (pixel_index <= 3794)) || ((pixel_index >= 3800) && (pixel_index <= 3801)) || ((pixel_index >= 3824) && (pixel_index <= 3833)) || ((pixel_index >= 3845) && (pixel_index <= 3871)) || ((pixel_index >= 3886) && (pixel_index <= 3890)) || pixel_index == 3896 || ((pixel_index >= 3921) && (pixel_index <= 3929)) || ((pixel_index >= 3941) && (pixel_index <= 3967)) || ((pixel_index >= 3982) && (pixel_index <= 3986)) || ((pixel_index >= 4017) && (pixel_index <= 4025)) || ((pixel_index >= 4037) && (pixel_index <= 4063)) || ((pixel_index >= 4078) && (pixel_index <= 4083)) || pixel_index == 4087 || pixel_index == 4111 || ((pixel_index >= 4113) && (pixel_index <= 4121)) || ((pixel_index >= 4133) && (pixel_index <= 4159)) || ((pixel_index >= 4174) && (pixel_index <= 4179)) || pixel_index == 4203 || pixel_index == 4205 || ((pixel_index >= 4207) && (pixel_index <= 4217)) || ((pixel_index >= 4229) && (pixel_index <= 4256)) || ((pixel_index >= 4270) && (pixel_index <= 4276)) || ((pixel_index >= 4299) && (pixel_index <= 4313)) || ((pixel_index >= 4325) && (pixel_index <= 4352)) || ((pixel_index >= 4367) && (pixel_index <= 4372)) || ((pixel_index >= 4395) && (pixel_index <= 4409)) || ((pixel_index >= 4421) && (pixel_index <= 4448)) || ((pixel_index >= 4464) && (pixel_index <= 4468)) || ((pixel_index >= 4492) && (pixel_index <= 4505)) || ((pixel_index >= 4517) && (pixel_index <= 4545)) || ((pixel_index >= 4561) && (pixel_index <= 4564)) || ((pixel_index >= 4588) && (pixel_index <= 4601)) || ((pixel_index >= 4613) && (pixel_index <= 4642)) || ((pixel_index >= 4658) && (pixel_index <= 4660)) || ((pixel_index >= 4684) && (pixel_index <= 4697)) || ((pixel_index >= 4709) && (pixel_index <= 4739)) || ((pixel_index >= 4781) && (pixel_index <= 4793)) || ((pixel_index >= 4805) && (pixel_index <= 4837)) || ((pixel_index >= 4878) && (pixel_index <= 4889)) || ((pixel_index >= 4901) && (pixel_index <= 4933)) || pixel_index == 4971 || ((pixel_index >= 4974) && (pixel_index <= 4985)) || ((pixel_index >= 4997) && (pixel_index <= 5029)) || ((pixel_index >= 5067) && (pixel_index <= 5081)) || ((pixel_index >= 5093) && (pixel_index <= 5124)) || ((pixel_index >= 5163) && (pixel_index <= 5177)) || ((pixel_index >= 5189) && (pixel_index <= 5220)) || ((pixel_index >= 5260) && (pixel_index <= 5273)) || ((pixel_index >= 5285) && (pixel_index <= 5316)) || ((pixel_index >= 5356) && (pixel_index <= 5369)) || ((pixel_index >= 5381) && (pixel_index <= 5412)) || ((pixel_index >= 5452) && (pixel_index <= 5465)) || ((pixel_index >= 5477) && (pixel_index <= 5507)) || ((pixel_index >= 5548) && (pixel_index <= 5561)) || ((pixel_index >= 5573) && (pixel_index <= 5603)) || ((pixel_index >= 5645) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5699)) || ((pixel_index >= 5741) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5795)) || ((pixel_index >= 5837) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5891)) || ((pixel_index >= 5933) && (pixel_index <= 5937)) || ((pixel_index >= 5941) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 5987)) || ((pixel_index >= 6029) && (pixel_index <= 6031)) || ((pixel_index >= 6036) && (pixel_index <= 6041)) || ((pixel_index >= 6053) && (pixel_index <= 6083)) || pixel_index == 6126 || (pixel_index >= 6132) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 11) begin
            if (((pixel_index >= 5) && (pixel_index <= 43)) || ((pixel_index >= 57) && (pixel_index <= 62)) || ((pixel_index >= 67) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 139)) || ((pixel_index >= 165) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 236)) || ((pixel_index >= 262) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 332)) || ((pixel_index >= 359) && (pixel_index <= 377)) || ((pixel_index >= 389) && (pixel_index <= 429)) || ((pixel_index >= 456) && (pixel_index <= 473)) || ((pixel_index >= 485) && (pixel_index <= 525)) || ((pixel_index >= 553) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 623)) || ((pixel_index >= 649) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 719)) || ((pixel_index >= 745) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 814)) || ((pixel_index >= 841) && (pixel_index <= 857)) || ((pixel_index >= 869) && (pixel_index <= 909)) || ((pixel_index >= 938) && (pixel_index <= 953)) || ((pixel_index >= 965) && (pixel_index <= 1004)) || ((pixel_index >= 1034) && (pixel_index <= 1049)) || ((pixel_index >= 1061) && (pixel_index <= 1099)) || ((pixel_index >= 1131) && (pixel_index <= 1145)) || ((pixel_index >= 1157) && (pixel_index <= 1194)) || ((pixel_index >= 1228) && (pixel_index <= 1241)) || ((pixel_index >= 1253) && (pixel_index <= 1290)) || ((pixel_index >= 1324) && (pixel_index <= 1337)) || ((pixel_index >= 1349) && (pixel_index <= 1385)) || ((pixel_index >= 1420) && (pixel_index <= 1433)) || ((pixel_index >= 1445) && (pixel_index <= 1481)) || ((pixel_index >= 1517) && (pixel_index <= 1529)) || ((pixel_index >= 1541) && (pixel_index <= 1577)) || ((pixel_index >= 1613) && (pixel_index <= 1625)) || ((pixel_index >= 1637) && (pixel_index <= 1673)) || ((pixel_index >= 1709) && (pixel_index <= 1721)) || ((pixel_index >= 1733) && (pixel_index <= 1768)) || ((pixel_index >= 1806) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1864)) || ((pixel_index >= 1902) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 1960)) || ((pixel_index >= 1998) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2056)) || ((pixel_index >= 2094) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2152)) || ((pixel_index >= 2190) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2248)) || ((pixel_index >= 2286) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2345)) || ((pixel_index >= 2382) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2442)) || ((pixel_index >= 2478) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2539)) || ((pixel_index >= 2574) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2636)) || ((pixel_index >= 2670) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2735)) || ((pixel_index >= 2766) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2832)) || ((pixel_index >= 2862) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2928)) || ((pixel_index >= 2958) && (pixel_index <= 2969)) || ((pixel_index >= 2981) && (pixel_index <= 3023)) || ((pixel_index >= 3054) && (pixel_index <= 3065)) || ((pixel_index >= 3077) && (pixel_index <= 3119)) || ((pixel_index >= 3150) && (pixel_index <= 3161)) || ((pixel_index >= 3173) && (pixel_index <= 3217)) || ((pixel_index >= 3246) && (pixel_index <= 3257)) || ((pixel_index >= 3269) && (pixel_index <= 3313)) || ((pixel_index >= 3342) && (pixel_index <= 3353)) || ((pixel_index >= 3365) && (pixel_index <= 3409)) || ((pixel_index >= 3438) && (pixel_index <= 3449)) || ((pixel_index >= 3461) && (pixel_index <= 3505)) || ((pixel_index >= 3513) && (pixel_index <= 3514)) || ((pixel_index >= 3534) && (pixel_index <= 3545)) || ((pixel_index >= 3557) && (pixel_index <= 3601)) || ((pixel_index >= 3608) && (pixel_index <= 3611)) || ((pixel_index >= 3630) && (pixel_index <= 3641)) || ((pixel_index >= 3653) && (pixel_index <= 3697)) || ((pixel_index >= 3704) && (pixel_index <= 3707)) || ((pixel_index >= 3726) && (pixel_index <= 3737)) || ((pixel_index >= 3749) && (pixel_index <= 3793)) || ((pixel_index >= 3799) && (pixel_index <= 3802)) || ((pixel_index >= 3823) && (pixel_index <= 3833)) || ((pixel_index >= 3845) && (pixel_index <= 3872)) || ((pixel_index >= 3880) && (pixel_index <= 3889)) || ((pixel_index >= 3895) && (pixel_index <= 3897)) || pixel_index == 3914 || ((pixel_index >= 3919) && (pixel_index <= 3929)) || ((pixel_index >= 3941) && (pixel_index <= 3967)) || ((pixel_index >= 3977) && (pixel_index <= 3985)) || ((pixel_index >= 3991) && (pixel_index <= 3993)) || pixel_index == 4010 || ((pixel_index >= 4015) && (pixel_index <= 4025)) || ((pixel_index >= 4037) && (pixel_index <= 4062)) || ((pixel_index >= 4073) && (pixel_index <= 4081)) || ((pixel_index >= 4087) && (pixel_index <= 4088)) || ((pixel_index >= 4106) && (pixel_index <= 4107)) || ((pixel_index >= 4110) && (pixel_index <= 4121)) || ((pixel_index >= 4133) && (pixel_index <= 4157)) || ((pixel_index >= 4170) && (pixel_index <= 4178)) || ((pixel_index >= 4182) && (pixel_index <= 4183)) || ((pixel_index >= 4202) && (pixel_index <= 4217)) || ((pixel_index >= 4229) && (pixel_index <= 4253)) || ((pixel_index >= 4266) && (pixel_index <= 4274)) || ((pixel_index >= 4278) && (pixel_index <= 4279)) || ((pixel_index >= 4299) && (pixel_index <= 4313)) || ((pixel_index >= 4325) && (pixel_index <= 4348)) || ((pixel_index >= 4362) && (pixel_index <= 4370)) || pixel_index == 4374 || ((pixel_index >= 4395) && (pixel_index <= 4409)) || ((pixel_index >= 4421) && (pixel_index <= 4444)) || ((pixel_index >= 4458) && (pixel_index <= 4466)) || pixel_index == 4470 || ((pixel_index >= 4491) && (pixel_index <= 4505)) || ((pixel_index >= 4517) && (pixel_index <= 4540)) || ((pixel_index >= 4555) && (pixel_index <= 4562)) || pixel_index == 4565 || ((pixel_index >= 4588) && (pixel_index <= 4601)) || ((pixel_index >= 4613) && (pixel_index <= 4636)) || ((pixel_index >= 4652) && (pixel_index <= 4658)) || pixel_index == 4661 || ((pixel_index >= 4684) && (pixel_index <= 4697)) || ((pixel_index >= 4709) && (pixel_index <= 4733)) || ((pixel_index >= 4749) && (pixel_index <= 4754)) || ((pixel_index >= 4778) && (pixel_index <= 4779)) || ((pixel_index >= 4781) && (pixel_index <= 4793)) || ((pixel_index >= 4805) && (pixel_index <= 4829)) || ((pixel_index >= 4847) && (pixel_index <= 4849)) || ((pixel_index >= 4874) && (pixel_index <= 4875)) || ((pixel_index >= 4878) && (pixel_index <= 4889)) || ((pixel_index >= 4901) && (pixel_index <= 4925)) || ((pixel_index >= 4944) && (pixel_index <= 4945)) || ((pixel_index >= 4970) && (pixel_index <= 4971)) || ((pixel_index >= 4974) && (pixel_index <= 4985)) || ((pixel_index >= 4997) && (pixel_index <= 5022)) || pixel_index == 5041 || ((pixel_index >= 5066) && (pixel_index <= 5068)) || ((pixel_index >= 5070) && (pixel_index <= 5081)) || ((pixel_index >= 5093) && (pixel_index <= 5119)) || ((pixel_index >= 5137) && (pixel_index <= 5138)) || ((pixel_index >= 5162) && (pixel_index <= 5177)) || ((pixel_index >= 5189) && (pixel_index <= 5216)) || ((pixel_index >= 5258) && (pixel_index <= 5273)) || ((pixel_index >= 5285) && (pixel_index <= 5314)) || ((pixel_index >= 5355) && (pixel_index <= 5369)) || ((pixel_index >= 5381) && (pixel_index <= 5413)) || ((pixel_index >= 5451) && (pixel_index <= 5465)) || ((pixel_index >= 5477) && (pixel_index <= 5508)) || ((pixel_index >= 5547) && (pixel_index <= 5561)) || ((pixel_index >= 5573) && (pixel_index <= 5604)) || ((pixel_index >= 5643) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5700)) || ((pixel_index >= 5739) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5795)) || ((pixel_index >= 5835) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5891)) || ((pixel_index >= 5932) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 5987)) || ((pixel_index >= 6028) && (pixel_index <= 6041)) || ((pixel_index >= 6053) && (pixel_index <= 6083)) || (pixel_index >= 6124) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 12) begin
            if (((pixel_index >= 5) && (pixel_index <= 34)) || ((pixel_index >= 49) && (pixel_index <= 50)) || ((pixel_index >= 65) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 130)) || ((pixel_index >= 162) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 226)) || ((pixel_index >= 259) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 323)) || ((pixel_index >= 356) && (pixel_index <= 377)) || ((pixel_index >= 389) && (pixel_index <= 419)) || ((pixel_index >= 452) && (pixel_index <= 473)) || ((pixel_index >= 485) && (pixel_index <= 516)) || ((pixel_index >= 549) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 613)) || ((pixel_index >= 646) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 710)) || ((pixel_index >= 743) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 807)) || ((pixel_index >= 839) && (pixel_index <= 857)) || ((pixel_index >= 869) && (pixel_index <= 904)) || ((pixel_index >= 936) && (pixel_index <= 953)) || ((pixel_index >= 965) && (pixel_index <= 1000)) || ((pixel_index >= 1033) && (pixel_index <= 1049)) || ((pixel_index >= 1061) && (pixel_index <= 1095)) || ((pixel_index >= 1129) && (pixel_index <= 1145)) || ((pixel_index >= 1157) && (pixel_index <= 1190)) || ((pixel_index >= 1226) && (pixel_index <= 1241)) || ((pixel_index >= 1253) && (pixel_index <= 1286)) || ((pixel_index >= 1322) && (pixel_index <= 1337)) || ((pixel_index >= 1349) && (pixel_index <= 1382)) || ((pixel_index >= 1419) && (pixel_index <= 1433)) || ((pixel_index >= 1445) && (pixel_index <= 1477)) || ((pixel_index >= 1515) && (pixel_index <= 1529)) || ((pixel_index >= 1541) && (pixel_index <= 1573)) || ((pixel_index >= 1611) && (pixel_index <= 1625)) || ((pixel_index >= 1637) && (pixel_index <= 1669)) || ((pixel_index >= 1708) && (pixel_index <= 1721)) || ((pixel_index >= 1733) && (pixel_index <= 1765)) || ((pixel_index >= 1804) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1861)) || ((pixel_index >= 1900) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 1957)) || ((pixel_index >= 1996) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2053)) || ((pixel_index >= 2093) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2149)) || ((pixel_index >= 2189) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2245)) || ((pixel_index >= 2285) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2341)) || ((pixel_index >= 2381) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2437)) || ((pixel_index >= 2478) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2534)) || ((pixel_index >= 2574) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2631)) || ((pixel_index >= 2670) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2729)) || ((pixel_index >= 2766) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2830)) || ((pixel_index >= 2862) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2926)) || ((pixel_index >= 2958) && (pixel_index <= 2969)) || ((pixel_index >= 2981) && (pixel_index <= 3022)) || ((pixel_index >= 3054) && (pixel_index <= 3065)) || ((pixel_index >= 3077) && (pixel_index <= 3118)) || ((pixel_index >= 3150) && (pixel_index <= 3161)) || ((pixel_index >= 3173) && (pixel_index <= 3215)) || ((pixel_index >= 3245) && (pixel_index <= 3257)) || ((pixel_index >= 3269) && (pixel_index <= 3311)) || ((pixel_index >= 3341) && (pixel_index <= 3353)) || ((pixel_index >= 3365) && (pixel_index <= 3407)) || pixel_index == 3417 || ((pixel_index >= 3437) && (pixel_index <= 3449)) || ((pixel_index >= 3461) && (pixel_index <= 3503)) || ((pixel_index >= 3513) && (pixel_index <= 3514)) || ((pixel_index >= 3534) && (pixel_index <= 3545)) || ((pixel_index >= 3557) && (pixel_index <= 3599)) || ((pixel_index >= 3609) && (pixel_index <= 3610)) || pixel_index == 3626 || ((pixel_index >= 3630) && (pixel_index <= 3641)) || ((pixel_index >= 3653) && (pixel_index <= 3695)) || pixel_index == 3701 || ((pixel_index >= 3705) && (pixel_index <= 3706)) || pixel_index == 3722 || ((pixel_index >= 3726) && (pixel_index <= 3737)) || ((pixel_index >= 3749) && (pixel_index <= 3792)) || pixel_index == 3797 || ((pixel_index >= 3801) && (pixel_index <= 3802)) || ((pixel_index >= 3818) && (pixel_index <= 3819)) || ((pixel_index >= 3823) && (pixel_index <= 3833)) || ((pixel_index >= 3845) && (pixel_index <= 3888)) || pixel_index == 3893 || pixel_index == 3897 || ((pixel_index >= 3914) && (pixel_index <= 3916)) || ((pixel_index >= 3919) && (pixel_index <= 3929)) || ((pixel_index >= 3941) && (pixel_index <= 3984)) || ((pixel_index >= 3989) && (pixel_index <= 3990)) || ((pixel_index >= 4010) && (pixel_index <= 4025)) || ((pixel_index >= 4037) && (pixel_index <= 4080)) || pixel_index == 4086 || ((pixel_index >= 4106) && (pixel_index <= 4121)) || ((pixel_index >= 4133) && (pixel_index <= 4176)) || ((pixel_index >= 4181) && (pixel_index <= 4182)) || ((pixel_index >= 4202) && (pixel_index <= 4217)) || ((pixel_index >= 4229) && (pixel_index <= 4273)) || ((pixel_index >= 4277) && (pixel_index <= 4278)) || ((pixel_index >= 4299) && (pixel_index <= 4313)) || ((pixel_index >= 4325) && (pixel_index <= 4369)) || pixel_index == 4373 || ((pixel_index >= 4395) && (pixel_index <= 4409)) || ((pixel_index >= 4421) && (pixel_index <= 4465)) || ((pixel_index >= 4468) && (pixel_index <= 4469)) || ((pixel_index >= 4491) && (pixel_index <= 4505)) || ((pixel_index >= 4517) && (pixel_index <= 4562)) || ((pixel_index >= 4588) && (pixel_index <= 4601)) || ((pixel_index >= 4613) && (pixel_index <= 4658)) || pixel_index == 4660 || ((pixel_index >= 4685) && (pixel_index <= 4697)) || ((pixel_index >= 4709) && (pixel_index <= 4754)) || pixel_index == 4756 || ((pixel_index >= 4782) && (pixel_index <= 4793)) || ((pixel_index >= 4805) && (pixel_index <= 4850)) || ((pixel_index >= 4878) && (pixel_index <= 4889)) || ((pixel_index >= 4901) && (pixel_index <= 4921)) || ((pixel_index >= 4928) && (pixel_index <= 4946)) || ((pixel_index >= 4974) && (pixel_index <= 4985)) || ((pixel_index >= 4997) && (pixel_index <= 5015)) || ((pixel_index >= 5025) && (pixel_index <= 5043)) || ((pixel_index >= 5069) && (pixel_index <= 5081)) || ((pixel_index >= 5093) && (pixel_index <= 5110)) || ((pixel_index >= 5122) && (pixel_index <= 5139)) || ((pixel_index >= 5165) && (pixel_index <= 5177)) || ((pixel_index >= 5189) && (pixel_index <= 5205)) || ((pixel_index >= 5218) && (pixel_index <= 5234)) || ((pixel_index >= 5262) && (pixel_index <= 5273)) || ((pixel_index >= 5285) && (pixel_index <= 5301)) || ((pixel_index >= 5314) && (pixel_index <= 5330)) || ((pixel_index >= 5358) && (pixel_index <= 5369)) || ((pixel_index >= 5381) && (pixel_index <= 5396)) || ((pixel_index >= 5410) && (pixel_index <= 5426)) || ((pixel_index >= 5454) && (pixel_index <= 5465)) || ((pixel_index >= 5477) && (pixel_index <= 5492)) || ((pixel_index >= 5506) && (pixel_index <= 5522)) || ((pixel_index >= 5550) && (pixel_index <= 5561)) || ((pixel_index >= 5573) && (pixel_index <= 5588)) || ((pixel_index >= 5603) && (pixel_index <= 5618)) || ((pixel_index >= 5646) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5685)) || ((pixel_index >= 5700) && (pixel_index <= 5714)) || ((pixel_index >= 5743) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5781)) || ((pixel_index >= 5807) && (pixel_index <= 5809)) || ((pixel_index >= 5839) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5877)) || ((pixel_index >= 5935) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 5973)) || ((pixel_index >= 6031) && (pixel_index <= 6041)) || ((pixel_index >= 6053) && (pixel_index <= 6070)) || (pixel_index >= 6127) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 13) begin
            if (((pixel_index >= 5) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 150)) || ((pixel_index >= 156) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 244)) || ((pixel_index >= 254) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 339)) || ((pixel_index >= 352) && (pixel_index <= 377)) || ((pixel_index >= 389) && (pixel_index <= 417)) || ((pixel_index >= 429) && (pixel_index <= 431)) || ((pixel_index >= 449) && (pixel_index <= 473)) || ((pixel_index >= 485) && (pixel_index <= 512)) || ((pixel_index >= 546) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 607)) || ((pixel_index >= 643) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 702)) || ((pixel_index >= 739) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 798)) || ((pixel_index >= 835) && (pixel_index <= 857)) || ((pixel_index >= 869) && (pixel_index <= 895)) || ((pixel_index >= 932) && (pixel_index <= 953)) || ((pixel_index >= 965) && (pixel_index <= 992)) || ((pixel_index >= 1029) && (pixel_index <= 1049)) || ((pixel_index >= 1061) && (pixel_index <= 1088)) || ((pixel_index >= 1126) && (pixel_index <= 1145)) || ((pixel_index >= 1157) && (pixel_index <= 1185)) || ((pixel_index >= 1222) && (pixel_index <= 1241)) || ((pixel_index >= 1253) && (pixel_index <= 1282)) || ((pixel_index >= 1319) && (pixel_index <= 1337)) || ((pixel_index >= 1349) && (pixel_index <= 1380)) || ((pixel_index >= 1416) && (pixel_index <= 1433)) || ((pixel_index >= 1445) && (pixel_index <= 1477)) || ((pixel_index >= 1512) && (pixel_index <= 1529)) || ((pixel_index >= 1541) && (pixel_index <= 1574)) || ((pixel_index >= 1608) && (pixel_index <= 1625)) || ((pixel_index >= 1637) && (pixel_index <= 1669)) || ((pixel_index >= 1705) && (pixel_index <= 1721)) || ((pixel_index >= 1733) && (pixel_index <= 1765)) || ((pixel_index >= 1801) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1860)) || ((pixel_index >= 1898) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 1956)) || ((pixel_index >= 1994) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2052)) || ((pixel_index >= 2090) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2148)) || ((pixel_index >= 2187) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2244)) || ((pixel_index >= 2283) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2340)) || ((pixel_index >= 2379) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2436)) || ((pixel_index >= 2475) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2532)) || ((pixel_index >= 2572) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2629)) || ((pixel_index >= 2668) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2725)) || ((pixel_index >= 2764) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2821)) || ((pixel_index >= 2861) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2917)) || ((pixel_index >= 2957) && (pixel_index <= 2969)) || ((pixel_index >= 2981) && (pixel_index <= 3014)) || ((pixel_index >= 3053) && (pixel_index <= 3065)) || ((pixel_index >= 3077) && (pixel_index <= 3111)) || ((pixel_index >= 3149) && (pixel_index <= 3161)) || ((pixel_index >= 3173) && (pixel_index <= 3209)) || ((pixel_index >= 3246) && (pixel_index <= 3257)) || ((pixel_index >= 3269) && (pixel_index <= 3309)) || ((pixel_index >= 3342) && (pixel_index <= 3353)) || ((pixel_index >= 3365) && (pixel_index <= 3405)) || ((pixel_index >= 3438) && (pixel_index <= 3449)) || ((pixel_index >= 3461) && (pixel_index <= 3501)) || ((pixel_index >= 3534) && (pixel_index <= 3545)) || ((pixel_index >= 3557) && (pixel_index <= 3597)) || ((pixel_index >= 3631) && (pixel_index <= 3641)) || ((pixel_index >= 3653) && (pixel_index <= 3693)) || pixel_index == 3697 || ((pixel_index >= 3725) && (pixel_index <= 3737)) || ((pixel_index >= 3749) && (pixel_index <= 3788)) || ((pixel_index >= 3793) && (pixel_index <= 3795)) || ((pixel_index >= 3801) && (pixel_index <= 3802)) || ((pixel_index >= 3822) && (pixel_index <= 3833)) || ((pixel_index >= 3845) && (pixel_index <= 3884)) || ((pixel_index >= 3890) && (pixel_index <= 3891)) || ((pixel_index >= 3896) && (pixel_index <= 3898)) || ((pixel_index >= 3917) && (pixel_index <= 3929)) || ((pixel_index >= 3941) && (pixel_index <= 3980)) || ((pixel_index >= 3985) && (pixel_index <= 3987)) || ((pixel_index >= 3991) && (pixel_index <= 3994)) || ((pixel_index >= 4013) && (pixel_index <= 4025)) || ((pixel_index >= 4037) && (pixel_index <= 4076)) || ((pixel_index >= 4081) && (pixel_index <= 4083)) || ((pixel_index >= 4088) && (pixel_index <= 4091)) || ((pixel_index >= 4110) && (pixel_index <= 4121)) || ((pixel_index >= 4133) && (pixel_index <= 4172)) || ((pixel_index >= 4177) && (pixel_index <= 4180)) || ((pixel_index >= 4183) && (pixel_index <= 4187)) || ((pixel_index >= 4206) && (pixel_index <= 4217)) || ((pixel_index >= 4229) && (pixel_index <= 4268)) || ((pixel_index >= 4273) && (pixel_index <= 4276)) || ((pixel_index >= 4279) && (pixel_index <= 4283)) || pixel_index == 4301 || ((pixel_index >= 4303) && (pixel_index <= 4313)) || ((pixel_index >= 4325) && (pixel_index <= 4364)) || ((pixel_index >= 4369) && (pixel_index <= 4373)) || ((pixel_index >= 4375) && (pixel_index <= 4378)) || ((pixel_index >= 4397) && (pixel_index <= 4409)) || ((pixel_index >= 4421) && (pixel_index <= 4460)) || ((pixel_index >= 4465) && (pixel_index <= 4469)) || ((pixel_index >= 4471) && (pixel_index <= 4473)) || ((pixel_index >= 4494) && (pixel_index <= 4505)) || ((pixel_index >= 4517) && (pixel_index <= 4556)) || ((pixel_index >= 4561) && (pixel_index <= 4565)) || ((pixel_index >= 4567) && (pixel_index <= 4569)) || ((pixel_index >= 4590) && (pixel_index <= 4601)) || ((pixel_index >= 4613) && (pixel_index <= 4652)) || ((pixel_index >= 4657) && (pixel_index <= 4664)) || ((pixel_index >= 4687) && (pixel_index <= 4697)) || ((pixel_index >= 4709) && (pixel_index <= 4749)) || ((pixel_index >= 4753) && (pixel_index <= 4760)) || ((pixel_index >= 4783) && (pixel_index <= 4793)) || ((pixel_index >= 4805) && (pixel_index <= 4845)) || ((pixel_index >= 4849) && (pixel_index <= 4855)) || ((pixel_index >= 4880) && (pixel_index <= 4889)) || ((pixel_index >= 4901) && (pixel_index <= 4942)) || ((pixel_index >= 4945) && (pixel_index <= 4950)) || ((pixel_index >= 4977) && (pixel_index <= 4985)) || ((pixel_index >= 4997) && (pixel_index <= 5038)) || ((pixel_index >= 5041) && (pixel_index <= 5046)) || ((pixel_index >= 5073) && (pixel_index <= 5081)) || ((pixel_index >= 5093) && (pixel_index <= 5134)) || ((pixel_index >= 5137) && (pixel_index <= 5141)) || ((pixel_index >= 5170) && (pixel_index <= 5177)) || ((pixel_index >= 5189) && (pixel_index <= 5231)) || ((pixel_index >= 5233) && (pixel_index <= 5237)) || ((pixel_index >= 5266) && (pixel_index <= 5273)) || ((pixel_index >= 5285) && (pixel_index <= 5327)) || ((pixel_index >= 5329) && (pixel_index <= 5333)) || ((pixel_index >= 5363) && (pixel_index <= 5369)) || ((pixel_index >= 5381) && (pixel_index <= 5429)) || ((pixel_index >= 5459) && (pixel_index <= 5465)) || ((pixel_index >= 5477) && (pixel_index <= 5525)) || ((pixel_index >= 5556) && (pixel_index <= 5561)) || ((pixel_index >= 5573) && (pixel_index <= 5621)) || ((pixel_index >= 5653) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5717)) || ((pixel_index >= 5749) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5813)) || ((pixel_index >= 5846) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5909)) || ((pixel_index >= 5942) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 6005)) || ((pixel_index >= 6039) && (pixel_index <= 6041)) || ((pixel_index >= 6053) && (pixel_index <= 6101)) || (pixel_index >= 6135) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 14) begin
            if (((pixel_index >= 5) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 377)) || ((pixel_index >= 389) && (pixel_index <= 473)) || ((pixel_index >= 485) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 821)) || ((pixel_index >= 828) && (pixel_index <= 857)) || ((pixel_index >= 869) && (pixel_index <= 916)) || ((pixel_index >= 926) && (pixel_index <= 927)) || ((pixel_index >= 930) && (pixel_index <= 932)) || ((pixel_index >= 939) && (pixel_index <= 953)) || ((pixel_index >= 965) && (pixel_index <= 1010)) || ((pixel_index >= 1037) && (pixel_index <= 1049)) || ((pixel_index >= 1061) && (pixel_index <= 1106)) || ((pixel_index >= 1134) && (pixel_index <= 1145)) || ((pixel_index >= 1157) && (pixel_index <= 1202)) || ((pixel_index >= 1231) && (pixel_index <= 1241)) || ((pixel_index >= 1253) && (pixel_index <= 1298)) || ((pixel_index >= 1327) && (pixel_index <= 1337)) || ((pixel_index >= 1349) && (pixel_index <= 1394)) || ((pixel_index >= 1424) && (pixel_index <= 1433)) || ((pixel_index >= 1445) && (pixel_index <= 1490)) || ((pixel_index >= 1521) && (pixel_index <= 1529)) || ((pixel_index >= 1541) && (pixel_index <= 1587)) || ((pixel_index >= 1617) && (pixel_index <= 1625)) || ((pixel_index >= 1637) && (pixel_index <= 1683)) || ((pixel_index >= 1713) && (pixel_index <= 1721)) || ((pixel_index >= 1733) && (pixel_index <= 1778)) || ((pixel_index >= 1809) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1873)) || ((pixel_index >= 1905) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 1968)) || ((pixel_index >= 2002) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2063)) || ((pixel_index >= 2098) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2159)) || ((pixel_index >= 2195) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2255)) || ((pixel_index >= 2291) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2350)) || ((pixel_index >= 2387) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2446)) || ((pixel_index >= 2483) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2542)) || ((pixel_index >= 2580) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2638)) || ((pixel_index >= 2676) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2734)) || ((pixel_index >= 2772) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2829)) || ((pixel_index >= 2868) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2925)) || ((pixel_index >= 2964) && (pixel_index <= 2969)) || ((pixel_index >= 2981) && (pixel_index <= 3021)) || ((pixel_index >= 3060) && (pixel_index <= 3065)) || ((pixel_index >= 3077) && (pixel_index <= 3118)) || ((pixel_index >= 3156) && (pixel_index <= 3161)) || ((pixel_index >= 3173) && (pixel_index <= 3214)) || ((pixel_index >= 3252) && (pixel_index <= 3257)) || ((pixel_index >= 3269) && (pixel_index <= 3311)) || ((pixel_index >= 3348) && (pixel_index <= 3353)) || ((pixel_index >= 3365) && (pixel_index <= 3408)) || ((pixel_index >= 3444) && (pixel_index <= 3449)) || ((pixel_index >= 3461) && (pixel_index <= 3506)) || ((pixel_index >= 3540) && (pixel_index <= 3545)) || ((pixel_index >= 3557) && (pixel_index <= 3604)) || ((pixel_index >= 3636) && (pixel_index <= 3641)) || ((pixel_index >= 3653) && (pixel_index <= 3701)) || ((pixel_index >= 3732) && (pixel_index <= 3737)) || ((pixel_index >= 3749) && (pixel_index <= 3797)) || ((pixel_index >= 3828) && (pixel_index <= 3833)) || ((pixel_index >= 3845) && (pixel_index <= 3892)) || ((pixel_index >= 3924) && (pixel_index <= 3929)) || ((pixel_index >= 3941) && (pixel_index <= 3989)) || ((pixel_index >= 4020) && (pixel_index <= 4025)) || ((pixel_index >= 4037) && (pixel_index <= 4085)) || ((pixel_index >= 4116) && (pixel_index <= 4121)) || ((pixel_index >= 4133) && (pixel_index <= 4180)) || ((pixel_index >= 4212) && (pixel_index <= 4217)) || ((pixel_index >= 4229) && (pixel_index <= 4275)) || ((pixel_index >= 4307) && (pixel_index <= 4313)) || ((pixel_index >= 4325) && (pixel_index <= 4371)) || ((pixel_index >= 4382) && (pixel_index <= 4383)) || ((pixel_index >= 4403) && (pixel_index <= 4409)) || ((pixel_index >= 4421) && (pixel_index <= 4466)) || pixel_index == 4474 || ((pixel_index >= 4476) && (pixel_index <= 4479)) || ((pixel_index >= 4499) && (pixel_index <= 4505)) || ((pixel_index >= 4517) && (pixel_index <= 4562)) || ((pixel_index >= 4570) && (pixel_index <= 4576)) || ((pixel_index >= 4596) && (pixel_index <= 4601)) || ((pixel_index >= 4613) && (pixel_index <= 4658)) || ((pixel_index >= 4665) && (pixel_index <= 4672)) || ((pixel_index >= 4692) && (pixel_index <= 4697)) || ((pixel_index >= 4709) && (pixel_index <= 4753)) || ((pixel_index >= 4760) && (pixel_index <= 4768)) || ((pixel_index >= 4789) && (pixel_index <= 4793)) || ((pixel_index >= 4805) && (pixel_index <= 4849)) || ((pixel_index >= 4856) && (pixel_index <= 4865)) || ((pixel_index >= 4886) && (pixel_index <= 4889)) || ((pixel_index >= 4901) && (pixel_index <= 4944)) || ((pixel_index >= 4952) && (pixel_index <= 4961)) || ((pixel_index >= 4982) && (pixel_index <= 4985)) || ((pixel_index >= 4997) && (pixel_index <= 5040)) || ((pixel_index >= 5047) && (pixel_index <= 5057)) || ((pixel_index >= 5079) && (pixel_index <= 5081)) || ((pixel_index >= 5093) && (pixel_index <= 5137)) || ((pixel_index >= 5143) && (pixel_index <= 5153)) || ((pixel_index >= 5176) && (pixel_index <= 5177)) || ((pixel_index >= 5189) && (pixel_index <= 5232)) || ((pixel_index >= 5236) && (pixel_index <= 5249)) || pixel_index == 5273 || ((pixel_index >= 5285) && (pixel_index <= 5328)) || ((pixel_index >= 5332) && (pixel_index <= 5344)) || pixel_index == 5369 || ((pixel_index >= 5381) && (pixel_index <= 5424)) || ((pixel_index >= 5427) && (pixel_index <= 5439)) || ((pixel_index >= 5477) && (pixel_index <= 5520)) || ((pixel_index >= 5522) && (pixel_index <= 5535)) || ((pixel_index >= 5573) && (pixel_index <= 5615)) || ((pixel_index >= 5618) && (pixel_index <= 5631)) || ((pixel_index >= 5669) && (pixel_index <= 5711)) || ((pixel_index >= 5713) && (pixel_index <= 5726)) || ((pixel_index >= 5765) && (pixel_index <= 5823)) || ((pixel_index >= 5861) && (pixel_index <= 5918)) || ((pixel_index >= 5957) && (pixel_index <= 6014)) || (pixel_index >= 6053) && (pixel_index <= 6110)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 15) begin
            if (((pixel_index >= 5) && (pixel_index <= 80)) || pixel_index == 89 || ((pixel_index >= 101) && (pixel_index <= 176)) || ((pixel_index >= 197) && (pixel_index <= 272)) || ((pixel_index >= 293) && (pixel_index <= 368)) || ((pixel_index >= 389) && (pixel_index <= 464)) || ((pixel_index >= 485) && (pixel_index <= 559)) || ((pixel_index >= 581) && (pixel_index <= 649)) || ((pixel_index >= 677) && (pixel_index <= 743)) || ((pixel_index >= 773) && (pixel_index <= 837)) || ((pixel_index >= 869) && (pixel_index <= 931)) || ((pixel_index >= 965) && (pixel_index <= 1026)) || ((pixel_index >= 1061) && (pixel_index <= 1121)) || ((pixel_index >= 1157) && (pixel_index <= 1216)) || ((pixel_index >= 1253) && (pixel_index <= 1312)) || ((pixel_index >= 1349) && (pixel_index <= 1407)) || ((pixel_index >= 1445) && (pixel_index <= 1503)) || ((pixel_index >= 1541) && (pixel_index <= 1598)) || ((pixel_index >= 1637) && (pixel_index <= 1694)) || ((pixel_index >= 1733) && (pixel_index <= 1789)) || ((pixel_index >= 1829) && (pixel_index <= 1886)) || ((pixel_index >= 1925) && (pixel_index <= 1982)) || ((pixel_index >= 2021) && (pixel_index <= 2078)) || ((pixel_index >= 2117) && (pixel_index <= 2174)) || ((pixel_index >= 2213) && (pixel_index <= 2270)) || ((pixel_index >= 2309) && (pixel_index <= 2367)) || ((pixel_index >= 2405) && (pixel_index <= 2464)) || ((pixel_index >= 2501) && (pixel_index <= 2562)) || ((pixel_index >= 2597) && (pixel_index <= 2658)) || ((pixel_index >= 2693) && (pixel_index <= 2753)) || ((pixel_index >= 2789) && (pixel_index <= 2848)) || ((pixel_index >= 2885) && (pixel_index <= 2945)) || ((pixel_index >= 2981) && (pixel_index <= 3042)) || ((pixel_index >= 3077) && (pixel_index <= 3138)) || ((pixel_index >= 3173) && (pixel_index <= 3235)) || ((pixel_index >= 3269) && (pixel_index <= 3331)) || ((pixel_index >= 3365) && (pixel_index <= 3427)) || ((pixel_index >= 3461) && (pixel_index <= 3523)) || ((pixel_index >= 3557) && (pixel_index <= 3619)) || pixel_index == 3624 || ((pixel_index >= 3653) && (pixel_index <= 3715)) || ((pixel_index >= 3719) && (pixel_index <= 3720)) || ((pixel_index >= 3749) && (pixel_index <= 3810)) || ((pixel_index >= 3815) && (pixel_index <= 3816)) || ((pixel_index >= 3845) && (pixel_index <= 3907)) || pixel_index == 3911 || ((pixel_index >= 3941) && (pixel_index <= 4003)) || ((pixel_index >= 4006) && (pixel_index <= 4008)) || ((pixel_index >= 4037) && (pixel_index <= 4099)) || ((pixel_index >= 4101) && (pixel_index <= 4104)) || ((pixel_index >= 4133) && (pixel_index <= 4195)) || ((pixel_index >= 4197) && (pixel_index <= 4200)) || ((pixel_index >= 4229) && (pixel_index <= 4291)) || ((pixel_index >= 4293) && (pixel_index <= 4296)) || ((pixel_index >= 4325) && (pixel_index <= 4392)) || ((pixel_index >= 4421) && (pixel_index <= 4488)) || ((pixel_index >= 4517) && (pixel_index <= 4583)) || ((pixel_index >= 4613) && (pixel_index <= 4679)) || ((pixel_index >= 4709) && (pixel_index <= 4775)) || ((pixel_index >= 4805) && (pixel_index <= 4871)) || ((pixel_index >= 4901) && (pixel_index <= 4967)) || ((pixel_index >= 4997) && (pixel_index <= 5064)) || ((pixel_index >= 5093) && (pixel_index <= 5160)) || ((pixel_index >= 5189) && (pixel_index <= 5256)) || ((pixel_index >= 5285) && (pixel_index <= 5352)) || ((pixel_index >= 5381) && (pixel_index <= 5448)) || ((pixel_index >= 5477) && (pixel_index <= 5544)) || ((pixel_index >= 5573) && (pixel_index <= 5640)) || ((pixel_index >= 5669) && (pixel_index <= 5735)) || ((pixel_index >= 5765) && (pixel_index <= 5831)) || ((pixel_index >= 5861) && (pixel_index <= 5927)) || ((pixel_index >= 5957) && (pixel_index <= 6023)) || (pixel_index >= 6053) && (pixel_index <= 6119)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 16) begin
            if (((pixel_index >= 5) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 376)) || ((pixel_index >= 389) && (pixel_index <= 470)) || ((pixel_index >= 485) && (pixel_index <= 564)) || ((pixel_index >= 581) && (pixel_index <= 659)) || ((pixel_index >= 677) && (pixel_index <= 753)) || ((pixel_index >= 773) && (pixel_index <= 849)) || ((pixel_index >= 869) && (pixel_index <= 944)) || ((pixel_index >= 965) && (pixel_index <= 1039)) || ((pixel_index >= 1061) && (pixel_index <= 1135)) || ((pixel_index >= 1157) && (pixel_index <= 1231)) || ((pixel_index >= 1253) && (pixel_index <= 1327)) || ((pixel_index >= 1349) && (pixel_index <= 1423)) || ((pixel_index >= 1445) && (pixel_index <= 1519)) || ((pixel_index >= 1541) && (pixel_index <= 1615)) || ((pixel_index >= 1637) && (pixel_index <= 1711)) || ((pixel_index >= 1733) && (pixel_index <= 1807)) || ((pixel_index >= 1829) && (pixel_index <= 1902)) || ((pixel_index >= 1925) && (pixel_index <= 1997)) || ((pixel_index >= 2021) && (pixel_index <= 2094)) || ((pixel_index >= 2117) && (pixel_index <= 2189)) || ((pixel_index >= 2213) && (pixel_index <= 2285)) || ((pixel_index >= 2309) && (pixel_index <= 2381)) || ((pixel_index >= 2405) && (pixel_index <= 2477)) || ((pixel_index >= 2501) && (pixel_index <= 2573)) || ((pixel_index >= 2597) && (pixel_index <= 2669)) || ((pixel_index >= 2693) && (pixel_index <= 2766)) || ((pixel_index >= 2789) && (pixel_index <= 2864)) || ((pixel_index >= 2885) && (pixel_index <= 2901)) || ((pixel_index >= 2903) && (pixel_index <= 2962)) || ((pixel_index >= 2981) && (pixel_index <= 2996)) || ((pixel_index >= 3001) && (pixel_index <= 3058)) || ((pixel_index >= 3077) && (pixel_index <= 3090)) || ((pixel_index >= 3098) && (pixel_index <= 3154)) || ((pixel_index >= 3173) && (pixel_index <= 3185)) || ((pixel_index >= 3195) && (pixel_index <= 3249)) || ((pixel_index >= 3269) && (pixel_index <= 3281)) || ((pixel_index >= 3292) && (pixel_index <= 3330)) || ((pixel_index >= 3333) && (pixel_index <= 3340)) || ((pixel_index >= 3365) && (pixel_index <= 3376)) || ((pixel_index >= 3388) && (pixel_index <= 3425)) || ((pixel_index >= 3430) && (pixel_index <= 3434)) || ((pixel_index >= 3461) && (pixel_index <= 3472)) || ((pixel_index >= 3485) && (pixel_index <= 3491)) || ((pixel_index >= 3498) && (pixel_index <= 3521)) || ((pixel_index >= 3526) && (pixel_index <= 3530)) || ((pixel_index >= 3557) && (pixel_index <= 3567)) || ((pixel_index >= 3582) && (pixel_index <= 3586)) || ((pixel_index >= 3600) && (pixel_index <= 3615)) || ((pixel_index >= 3653) && (pixel_index <= 3663)) || ((pixel_index >= 3679) && (pixel_index <= 3681)) || ((pixel_index >= 3700) && (pixel_index <= 3706)) || ((pixel_index >= 3749) && (pixel_index <= 3759)) || ((pixel_index >= 3775) && (pixel_index <= 3776)) || ((pixel_index >= 3845) && (pixel_index <= 3855)) || ((pixel_index >= 3871) && (pixel_index <= 3872)) || ((pixel_index >= 3941) && (pixel_index <= 3952)) || ((pixel_index >= 3967) && (pixel_index <= 3968)) || ((pixel_index >= 4037) && (pixel_index <= 4048)) || ((pixel_index >= 4063) && (pixel_index <= 4064)) || ((pixel_index >= 4133) && (pixel_index <= 4145)) || ((pixel_index >= 4158) && (pixel_index <= 4160)) || ((pixel_index >= 4229) && (pixel_index <= 4242)) || ((pixel_index >= 4252) && (pixel_index <= 4257)) || ((pixel_index >= 4325) && (pixel_index <= 4353)) || ((pixel_index >= 4421) && (pixel_index <= 4449)) || pixel_index == 4481 || ((pixel_index >= 4517) && (pixel_index <= 4545)) || ((pixel_index >= 4575) && (pixel_index <= 4579)) || ((pixel_index >= 4613) && (pixel_index <= 4641)) || ((pixel_index >= 4670) && (pixel_index <= 4675)) || ((pixel_index >= 4709) && (pixel_index <= 4737)) || ((pixel_index >= 4766) && (pixel_index <= 4771)) || ((pixel_index >= 4805) && (pixel_index <= 4833)) || ((pixel_index >= 4862) && (pixel_index <= 4867)) || ((pixel_index >= 4901) && (pixel_index <= 4929)) || ((pixel_index >= 4958) && (pixel_index <= 4963)) || ((pixel_index >= 4997) && (pixel_index <= 5024)) || ((pixel_index >= 5055) && (pixel_index <= 5058)) || ((pixel_index >= 5093) && (pixel_index <= 5120)) || ((pixel_index >= 5151) && (pixel_index <= 5154)) || ((pixel_index >= 5189) && (pixel_index <= 5216)) || ((pixel_index >= 5247) && (pixel_index <= 5250)) || ((pixel_index >= 5285) && (pixel_index <= 5312)) || ((pixel_index >= 5344) && (pixel_index <= 5346)) || ((pixel_index >= 5381) && (pixel_index <= 5408)) || ((pixel_index >= 5440) && (pixel_index <= 5442)) || ((pixel_index >= 5477) && (pixel_index <= 5504)) || ((pixel_index >= 5537) && (pixel_index <= 5538)) || ((pixel_index >= 5573) && (pixel_index <= 5600)) || ((pixel_index >= 5633) && (pixel_index <= 5634)) || ((pixel_index >= 5669) && (pixel_index <= 5696)) || ((pixel_index >= 5729) && (pixel_index <= 5730)) || ((pixel_index >= 5765) && (pixel_index <= 5792)) || ((pixel_index >= 5825) && (pixel_index <= 5826)) || ((pixel_index >= 5861) && (pixel_index <= 5888)) || pixel_index == 5922 || ((pixel_index >= 5957) && (pixel_index <= 5984)) || pixel_index == 6018 || ((pixel_index >= 6053) && (pixel_index <= 6080)) || pixel_index == 6114) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 17) begin
            if (((pixel_index >= 5) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 377)) || ((pixel_index >= 389) && (pixel_index <= 473)) || ((pixel_index >= 485) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 857)) || ((pixel_index >= 869) && (pixel_index <= 953)) || ((pixel_index >= 965) && (pixel_index <= 1049)) || ((pixel_index >= 1061) && (pixel_index <= 1145)) || ((pixel_index >= 1157) && (pixel_index <= 1241)) || ((pixel_index >= 1253) && (pixel_index <= 1337)) || ((pixel_index >= 1349) && (pixel_index <= 1433)) || ((pixel_index >= 1445) && (pixel_index <= 1529)) || ((pixel_index >= 1541) && (pixel_index <= 1625)) || ((pixel_index >= 1637) && (pixel_index <= 1721)) || ((pixel_index >= 1733) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2969)) || ((pixel_index >= 2981) && (pixel_index <= 3065)) || ((pixel_index >= 3077) && (pixel_index <= 3146)) || ((pixel_index >= 3148) && (pixel_index <= 3161)) || ((pixel_index >= 3173) && (pixel_index <= 3240)) || ((pixel_index >= 3245) && (pixel_index <= 3257)) || ((pixel_index >= 3269) && (pixel_index <= 3326)) || ((pixel_index >= 3328) && (pixel_index <= 3336)) || ((pixel_index >= 3341) && (pixel_index <= 3353)) || ((pixel_index >= 3365) && (pixel_index <= 3421)) || ((pixel_index >= 3424) && (pixel_index <= 3432)) || ((pixel_index >= 3438) && (pixel_index <= 3449)) || ((pixel_index >= 3461) && (pixel_index <= 3517)) || ((pixel_index >= 3520) && (pixel_index <= 3527)) || ((pixel_index >= 3534) && (pixel_index <= 3545)) || ((pixel_index >= 3557) && (pixel_index <= 3613)) || ((pixel_index >= 3617) && (pixel_index <= 3623)) || ((pixel_index >= 3630) && (pixel_index <= 3641)) || ((pixel_index >= 3653) && (pixel_index <= 3709)) || ((pixel_index >= 3713) && (pixel_index <= 3718)) || ((pixel_index >= 3723) && (pixel_index <= 3724)) || ((pixel_index >= 3726) && (pixel_index <= 3737)) || ((pixel_index >= 3749) && (pixel_index <= 3804)) || ((pixel_index >= 3809) && (pixel_index <= 3814)) || ((pixel_index >= 3820) && (pixel_index <= 3833)) || ((pixel_index >= 3845) && (pixel_index <= 3900)) || ((pixel_index >= 3905) && (pixel_index <= 3909)) || ((pixel_index >= 3916) && (pixel_index <= 3929)) || ((pixel_index >= 3941) && (pixel_index <= 3996)) || ((pixel_index >= 4001) && (pixel_index <= 4005)) || ((pixel_index >= 4012) && (pixel_index <= 4025)) || ((pixel_index >= 4037) && (pixel_index <= 4092)) || ((pixel_index >= 4097) && (pixel_index <= 4100)) || ((pixel_index >= 4107) && (pixel_index <= 4121)) || ((pixel_index >= 4133) && (pixel_index <= 4187)) || ((pixel_index >= 4193) && (pixel_index <= 4196)) || ((pixel_index >= 4203) && (pixel_index <= 4217)) || ((pixel_index >= 4229) && (pixel_index <= 4283)) || ((pixel_index >= 4289) && (pixel_index <= 4291)) || ((pixel_index >= 4299) && (pixel_index <= 4313)) || ((pixel_index >= 4325) && (pixel_index <= 4378)) || ((pixel_index >= 4385) && (pixel_index <= 4387)) || ((pixel_index >= 4394) && (pixel_index <= 4409)) || ((pixel_index >= 4421) && (pixel_index <= 4473)) || ((pixel_index >= 4481) && (pixel_index <= 4482)) || ((pixel_index >= 4490) && (pixel_index <= 4505)) || ((pixel_index >= 4517) && (pixel_index <= 4569)) || ((pixel_index >= 4576) && (pixel_index <= 4578)) || ((pixel_index >= 4586) && (pixel_index <= 4601)) || ((pixel_index >= 4613) && (pixel_index <= 4664)) || pixel_index == 4673 || ((pixel_index >= 4682) && (pixel_index <= 4697)) || ((pixel_index >= 4709) && (pixel_index <= 4759)) || pixel_index == 4769 || ((pixel_index >= 4778) && (pixel_index <= 4793)) || ((pixel_index >= 4805) && (pixel_index <= 4855)) || ((pixel_index >= 4874) && (pixel_index <= 4889)) || ((pixel_index >= 4901) && (pixel_index <= 4950)) || ((pixel_index >= 4969) && (pixel_index <= 4985)) || ((pixel_index >= 4997) && (pixel_index <= 5045)) || ((pixel_index >= 5065) && (pixel_index <= 5081)) || ((pixel_index >= 5093) && (pixel_index <= 5140)) || ((pixel_index >= 5161) && (pixel_index <= 5177)) || ((pixel_index >= 5189) && (pixel_index <= 5235)) || ((pixel_index >= 5257) && (pixel_index <= 5273)) || ((pixel_index >= 5285) && (pixel_index <= 5331)) || ((pixel_index >= 5353) && (pixel_index <= 5369)) || ((pixel_index >= 5381) && (pixel_index <= 5426)) || ((pixel_index >= 5449) && (pixel_index <= 5465)) || ((pixel_index >= 5477) && (pixel_index <= 5522)) || ((pixel_index >= 5545) && (pixel_index <= 5561)) || ((pixel_index >= 5573) && (pixel_index <= 5617)) || ((pixel_index >= 5642) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5712)) || ((pixel_index >= 5738) && (pixel_index <= 5752)) || ((pixel_index >= 5765) && (pixel_index <= 5807)) || ((pixel_index >= 5834) && (pixel_index <= 5848)) || ((pixel_index >= 5861) && (pixel_index <= 5903)) || ((pixel_index >= 5930) && (pixel_index <= 5944)) || ((pixel_index >= 5957) && (pixel_index <= 5998)) || ((pixel_index >= 6026) && (pixel_index <= 6040)) || ((pixel_index >= 6053) && (pixel_index <= 6093)) || (pixel_index >= 6122) && (pixel_index <= 6136)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 18) begin
            if (((pixel_index >= 5) && (pixel_index <= 35)) || ((pixel_index >= 51) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 131)) || ((pixel_index >= 147) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 227)) || ((pixel_index >= 243) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 323)) || ((pixel_index >= 339) && (pixel_index <= 377)) || ((pixel_index >= 389) && (pixel_index <= 420)) || ((pixel_index >= 435) && (pixel_index <= 473)) || ((pixel_index >= 485) && (pixel_index <= 516)) || ((pixel_index >= 530) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 613)) || ((pixel_index >= 625) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 710)) || ((pixel_index >= 721) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 807)) || ((pixel_index >= 815) && (pixel_index <= 857)) || ((pixel_index >= 869) && (pixel_index <= 904)) || ((pixel_index >= 909) && (pixel_index <= 953)) || ((pixel_index >= 965) && (pixel_index <= 1049)) || ((pixel_index >= 1061) && (pixel_index <= 1145)) || ((pixel_index >= 1157) && (pixel_index <= 1241)) || ((pixel_index >= 1253) && (pixel_index <= 1337)) || ((pixel_index >= 1349) && (pixel_index <= 1433)) || ((pixel_index >= 1445) && (pixel_index <= 1529)) || ((pixel_index >= 1541) && (pixel_index <= 1625)) || ((pixel_index >= 1637) && (pixel_index <= 1721)) || ((pixel_index >= 1733) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2969)) || ((pixel_index >= 2981) && (pixel_index <= 3065)) || ((pixel_index >= 3077) && (pixel_index <= 3161)) || ((pixel_index >= 3173) && (pixel_index <= 3257)) || ((pixel_index >= 3269) && (pixel_index <= 3353)) || ((pixel_index >= 3365) && (pixel_index <= 3449)) || ((pixel_index >= 3461) && (pixel_index <= 3545)) || ((pixel_index >= 3557) && (pixel_index <= 3641)) || ((pixel_index >= 3653) && (pixel_index <= 3737)) || ((pixel_index >= 3749) && (pixel_index <= 3833)) || ((pixel_index >= 3845) && (pixel_index <= 3929)) || ((pixel_index >= 3941) && (pixel_index <= 4025)) || ((pixel_index >= 4037) && (pixel_index <= 4121)) || ((pixel_index >= 4133) && (pixel_index <= 4217)) || ((pixel_index >= 4229) && (pixel_index <= 4313)) || ((pixel_index >= 4325) && (pixel_index <= 4409)) || ((pixel_index >= 4421) && (pixel_index <= 4505)) || ((pixel_index >= 4517) && (pixel_index <= 4601)) || ((pixel_index >= 4613) && (pixel_index <= 4697)) || ((pixel_index >= 4709) && (pixel_index <= 4793)) || ((pixel_index >= 4805) && (pixel_index <= 4889)) || ((pixel_index >= 4901) && (pixel_index <= 4985)) || ((pixel_index >= 4997) && (pixel_index <= 5081)) || ((pixel_index >= 5093) && (pixel_index <= 5177)) || ((pixel_index >= 5189) && (pixel_index <= 5273)) || ((pixel_index >= 5285) && (pixel_index <= 5369)) || ((pixel_index >= 5381) && (pixel_index <= 5465)) || ((pixel_index >= 5477) && (pixel_index <= 5561)) || ((pixel_index >= 5573) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 6041)) || (pixel_index >= 6053) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 19) begin
            if (((pixel_index >= 5) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 377)) || ((pixel_index >= 389) && (pixel_index <= 473)) || ((pixel_index >= 485) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 813)) || ((pixel_index >= 816) && (pixel_index <= 857)) || ((pixel_index >= 869) && (pixel_index <= 907)) || ((pixel_index >= 915) && (pixel_index <= 953)) || ((pixel_index >= 965) && (pixel_index <= 1001)) || ((pixel_index >= 1013) && (pixel_index <= 1049)) || ((pixel_index >= 1061) && (pixel_index <= 1096)) || ((pixel_index >= 1110) && (pixel_index <= 1145)) || ((pixel_index >= 1157) && (pixel_index <= 1191)) || ((pixel_index >= 1207) && (pixel_index <= 1241)) || ((pixel_index >= 1253) && (pixel_index <= 1287)) || ((pixel_index >= 1303) && (pixel_index <= 1337)) || ((pixel_index >= 1349) && (pixel_index <= 1382)) || ((pixel_index >= 1400) && (pixel_index <= 1433)) || ((pixel_index >= 1445) && (pixel_index <= 1478)) || ((pixel_index >= 1496) && (pixel_index <= 1529)) || ((pixel_index >= 1541) && (pixel_index <= 1573)) || ((pixel_index >= 1592) && (pixel_index <= 1625)) || ((pixel_index >= 1637) && (pixel_index <= 1669)) || ((pixel_index >= 1689) && (pixel_index <= 1721)) || ((pixel_index >= 1733) && (pixel_index <= 1765)) || ((pixel_index >= 1785) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1861)) || ((pixel_index >= 1881) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 1957)) || ((pixel_index >= 1976) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2054)) || ((pixel_index >= 2072) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2150)) || ((pixel_index >= 2167) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2247)) || ((pixel_index >= 2262) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2343)) || ((pixel_index >= 2357) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2441)) || ((pixel_index >= 2452) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2538)) || ((pixel_index >= 2546) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2969)) || ((pixel_index >= 2981) && (pixel_index <= 3065)) || ((pixel_index >= 3077) && (pixel_index <= 3161)) || ((pixel_index >= 3173) && (pixel_index <= 3257)) || ((pixel_index >= 3269) && (pixel_index <= 3353)) || ((pixel_index >= 3365) && (pixel_index <= 3449)) || ((pixel_index >= 3461) && (pixel_index <= 3545)) || ((pixel_index >= 3557) && (pixel_index <= 3641)) || ((pixel_index >= 3653) && (pixel_index <= 3737)) || ((pixel_index >= 3749) && (pixel_index <= 3833)) || ((pixel_index >= 3845) && (pixel_index <= 3929)) || ((pixel_index >= 3941) && (pixel_index <= 4025)) || ((pixel_index >= 4037) && (pixel_index <= 4121)) || ((pixel_index >= 4133) && (pixel_index <= 4217)) || ((pixel_index >= 4229) && (pixel_index <= 4313)) || ((pixel_index >= 4325) && (pixel_index <= 4409)) || ((pixel_index >= 4421) && (pixel_index <= 4505)) || ((pixel_index >= 4517) && (pixel_index <= 4601)) || ((pixel_index >= 4613) && (pixel_index <= 4697)) || ((pixel_index >= 4709) && (pixel_index <= 4793)) || ((pixel_index >= 4805) && (pixel_index <= 4889)) || ((pixel_index >= 4901) && (pixel_index <= 4985)) || ((pixel_index >= 4997) && (pixel_index <= 5081)) || ((pixel_index >= 5093) && (pixel_index <= 5177)) || ((pixel_index >= 5189) && (pixel_index <= 5273)) || ((pixel_index >= 5285) && (pixel_index <= 5369)) || ((pixel_index >= 5381) && (pixel_index <= 5465)) || ((pixel_index >= 5477) && (pixel_index <= 5561)) || ((pixel_index >= 5573) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 6041)) || (pixel_index >= 6053) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 20) begin
            if (((pixel_index >= 5) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 377)) || ((pixel_index >= 389) && (pixel_index <= 473)) || ((pixel_index >= 485) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 857)) || ((pixel_index >= 869) && (pixel_index <= 953)) || ((pixel_index >= 965) && (pixel_index <= 1049)) || ((pixel_index >= 1061) && (pixel_index <= 1145)) || ((pixel_index >= 1157) && (pixel_index <= 1241)) || ((pixel_index >= 1253) && (pixel_index <= 1337)) || ((pixel_index >= 1349) && (pixel_index <= 1433)) || ((pixel_index >= 1445) && (pixel_index <= 1529)) || ((pixel_index >= 1541) && (pixel_index <= 1625)) || ((pixel_index >= 1637) && (pixel_index <= 1721)) || ((pixel_index >= 1733) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2063)) || ((pixel_index >= 2068) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2157)) || ((pixel_index >= 2166) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2252)) || ((pixel_index >= 2263) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2348)) || ((pixel_index >= 2361) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2443)) || ((pixel_index >= 2457) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2535)) || ((pixel_index >= 2537) && (pixel_index <= 2538)) || ((pixel_index >= 2554) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2633)) || ((pixel_index >= 2651) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2729)) || ((pixel_index >= 2748) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2825)) || ((pixel_index >= 2844) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2920)) || ((pixel_index >= 2940) && (pixel_index <= 2969)) || ((pixel_index >= 2981) && (pixel_index <= 3016)) || ((pixel_index >= 3037) && (pixel_index <= 3065)) || ((pixel_index >= 3077) && (pixel_index <= 3111)) || ((pixel_index >= 3133) && (pixel_index <= 3161)) || ((pixel_index >= 3173) && (pixel_index <= 3207)) || ((pixel_index >= 3228) && (pixel_index <= 3257)) || ((pixel_index >= 3269) && (pixel_index <= 3304)) || ((pixel_index >= 3323) && (pixel_index <= 3353)) || ((pixel_index >= 3365) && (pixel_index <= 3400)) || ((pixel_index >= 3419) && (pixel_index <= 3449)) || ((pixel_index >= 3461) && (pixel_index <= 3496)) || ((pixel_index >= 3515) && (pixel_index <= 3545)) || ((pixel_index >= 3557) && (pixel_index <= 3593)) || ((pixel_index >= 3611) && (pixel_index <= 3641)) || ((pixel_index >= 3653) && (pixel_index <= 3689)) || ((pixel_index >= 3706) && (pixel_index <= 3737)) || ((pixel_index >= 3749) && (pixel_index <= 3787)) || ((pixel_index >= 3801) && (pixel_index <= 3833)) || ((pixel_index >= 3845) && (pixel_index <= 3885)) || ((pixel_index >= 3896) && (pixel_index <= 3929)) || ((pixel_index >= 3941) && (pixel_index <= 3984)) || ((pixel_index >= 3990) && (pixel_index <= 4025)) || ((pixel_index >= 4037) && (pixel_index <= 4121)) || ((pixel_index >= 4133) && (pixel_index <= 4217)) || ((pixel_index >= 4229) && (pixel_index <= 4313)) || ((pixel_index >= 4325) && (pixel_index <= 4409)) || ((pixel_index >= 4421) && (pixel_index <= 4505)) || ((pixel_index >= 4517) && (pixel_index <= 4601)) || ((pixel_index >= 4613) && (pixel_index <= 4697)) || ((pixel_index >= 4709) && (pixel_index <= 4793)) || ((pixel_index >= 4805) && (pixel_index <= 4889)) || ((pixel_index >= 4901) && (pixel_index <= 4985)) || ((pixel_index >= 4997) && (pixel_index <= 5081)) || ((pixel_index >= 5093) && (pixel_index <= 5177)) || ((pixel_index >= 5189) && (pixel_index <= 5273)) || ((pixel_index >= 5285) && (pixel_index <= 5369)) || ((pixel_index >= 5381) && (pixel_index <= 5465)) || ((pixel_index >= 5477) && (pixel_index <= 5561)) || ((pixel_index >= 5573) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 6041)) || (pixel_index >= 6053) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 21) begin
            if (((pixel_index >= 5) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 377)) || ((pixel_index >= 389) && (pixel_index <= 473)) || ((pixel_index >= 485) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 857)) || ((pixel_index >= 869) && (pixel_index <= 953)) || ((pixel_index >= 965) && (pixel_index <= 1049)) || ((pixel_index >= 1061) && (pixel_index <= 1145)) || ((pixel_index >= 1157) && (pixel_index <= 1241)) || ((pixel_index >= 1253) && (pixel_index <= 1337)) || ((pixel_index >= 1349) && (pixel_index <= 1433)) || ((pixel_index >= 1445) && (pixel_index <= 1529)) || ((pixel_index >= 1541) && (pixel_index <= 1625)) || ((pixel_index >= 1637) && (pixel_index <= 1721)) || ((pixel_index >= 1733) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2928)) || ((pixel_index >= 2933) && (pixel_index <= 2969)) || ((pixel_index >= 2981) && (pixel_index <= 3023)) || ((pixel_index >= 3032) && (pixel_index <= 3065)) || ((pixel_index >= 3077) && (pixel_index <= 3117)) || ((pixel_index >= 3130) && (pixel_index <= 3161)) || ((pixel_index >= 3173) && (pixel_index <= 3212)) || ((pixel_index >= 3227) && (pixel_index <= 3257)) || ((pixel_index >= 3269) && (pixel_index <= 3307)) || ((pixel_index >= 3324) && (pixel_index <= 3353)) || ((pixel_index >= 3365) && (pixel_index <= 3402)) || ((pixel_index >= 3421) && (pixel_index <= 3449)) || ((pixel_index >= 3461) && (pixel_index <= 3498)) || ((pixel_index >= 3517) && (pixel_index <= 3545)) || ((pixel_index >= 3557) && (pixel_index <= 3593)) || ((pixel_index >= 3613) && (pixel_index <= 3641)) || ((pixel_index >= 3653) && (pixel_index <= 3689)) || ((pixel_index >= 3709) && (pixel_index <= 3737)) || ((pixel_index >= 3749) && (pixel_index <= 3785)) || ((pixel_index >= 3806) && (pixel_index <= 3833)) || ((pixel_index >= 3845) && (pixel_index <= 3880)) || ((pixel_index >= 3902) && (pixel_index <= 3929)) || ((pixel_index >= 3941) && (pixel_index <= 3976)) || ((pixel_index >= 3998) && (pixel_index <= 4025)) || ((pixel_index >= 4037) && (pixel_index <= 4072)) || ((pixel_index >= 4094) && (pixel_index <= 4121)) || ((pixel_index >= 4133) && (pixel_index <= 4168)) || ((pixel_index >= 4190) && (pixel_index <= 4217)) || ((pixel_index >= 4229) && (pixel_index <= 4264)) || ((pixel_index >= 4286) && (pixel_index <= 4313)) || ((pixel_index >= 4325) && (pixel_index <= 4360)) || ((pixel_index >= 4381) && (pixel_index <= 4409)) || ((pixel_index >= 4421) && (pixel_index <= 4457)) || ((pixel_index >= 4477) && (pixel_index <= 4505)) || ((pixel_index >= 4517) && (pixel_index <= 4554)) || ((pixel_index >= 4573) && (pixel_index <= 4601)) || ((pixel_index >= 4613) && (pixel_index <= 4651)) || ((pixel_index >= 4668) && (pixel_index <= 4697)) || ((pixel_index >= 4709) && (pixel_index <= 4749)) || ((pixel_index >= 4763) && (pixel_index <= 4793)) || ((pixel_index >= 4805) && (pixel_index <= 4847)) || ((pixel_index >= 4857) && (pixel_index <= 4889)) || ((pixel_index >= 4901) && (pixel_index <= 4944)) || ((pixel_index >= 4946) && (pixel_index <= 4985)) || ((pixel_index >= 4997) && (pixel_index <= 5081)) || ((pixel_index >= 5093) && (pixel_index <= 5135)) || ((pixel_index >= 5137) && (pixel_index <= 5177)) || ((pixel_index >= 5189) && (pixel_index <= 5273)) || ((pixel_index >= 5285) && (pixel_index <= 5369)) || ((pixel_index >= 5381) && (pixel_index <= 5465)) || ((pixel_index >= 5477) && (pixel_index <= 5561)) || ((pixel_index >= 5573) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 6041)) || (pixel_index >= 6053) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 22) begin
            if (((pixel_index >= 5) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 377)) || ((pixel_index >= 389) && (pixel_index <= 473)) || ((pixel_index >= 485) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 857)) || ((pixel_index >= 869) && (pixel_index <= 953)) || ((pixel_index >= 965) && (pixel_index <= 1049)) || ((pixel_index >= 1061) && (pixel_index <= 1145)) || ((pixel_index >= 1157) && (pixel_index <= 1241)) || ((pixel_index >= 1253) && (pixel_index <= 1337)) || ((pixel_index >= 1349) && (pixel_index <= 1433)) || ((pixel_index >= 1445) && (pixel_index <= 1529)) || ((pixel_index >= 1541) && (pixel_index <= 1625)) || ((pixel_index >= 1637) && (pixel_index <= 1721)) || ((pixel_index >= 1733) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2969)) || ((pixel_index >= 2981) && (pixel_index <= 3065)) || ((pixel_index >= 3077) && (pixel_index <= 3161)) || ((pixel_index >= 3173) && (pixel_index <= 3257)) || ((pixel_index >= 3269) && (pixel_index <= 3353)) || ((pixel_index >= 3365) && (pixel_index <= 3407)) || ((pixel_index >= 3418) && (pixel_index <= 3449)) || ((pixel_index >= 3461) && (pixel_index <= 3501)) || ((pixel_index >= 3515) && (pixel_index <= 3545)) || ((pixel_index >= 3557) && (pixel_index <= 3595)) || ((pixel_index >= 3612) && (pixel_index <= 3641)) || ((pixel_index >= 3653) && (pixel_index <= 3690)) || ((pixel_index >= 3709) && (pixel_index <= 3737)) || ((pixel_index >= 3749) && (pixel_index <= 3785)) || ((pixel_index >= 3805) && (pixel_index <= 3833)) || ((pixel_index >= 3845) && (pixel_index <= 3881)) || ((pixel_index >= 3902) && (pixel_index <= 3929)) || ((pixel_index >= 3941) && (pixel_index <= 3977)) || ((pixel_index >= 3998) && (pixel_index <= 4025)) || ((pixel_index >= 4037) && (pixel_index <= 4073)) || ((pixel_index >= 4094) && (pixel_index <= 4121)) || ((pixel_index >= 4133) && (pixel_index <= 4168)) || ((pixel_index >= 4190) && (pixel_index <= 4217)) || ((pixel_index >= 4229) && (pixel_index <= 4265)) || ((pixel_index >= 4286) && (pixel_index <= 4313)) || ((pixel_index >= 4325) && (pixel_index <= 4361)) || ((pixel_index >= 4383) && (pixel_index <= 4409)) || ((pixel_index >= 4421) && (pixel_index <= 4456)) || ((pixel_index >= 4480) && (pixel_index <= 4505)) || ((pixel_index >= 4517) && (pixel_index <= 4552)) || ((pixel_index >= 4574) && (pixel_index <= 4601)) || ((pixel_index >= 4613) && (pixel_index <= 4648)) || ((pixel_index >= 4670) && (pixel_index <= 4697)) || ((pixel_index >= 4709) && (pixel_index <= 4744)) || ((pixel_index >= 4765) && (pixel_index <= 4793)) || ((pixel_index >= 4805) && (pixel_index <= 4841)) || ((pixel_index >= 4861) && (pixel_index <= 4889)) || ((pixel_index >= 4901) && (pixel_index <= 4938)) || ((pixel_index >= 4957) && (pixel_index <= 4985)) || ((pixel_index >= 4997) && (pixel_index <= 5035)) || ((pixel_index >= 5053) && (pixel_index <= 5081)) || ((pixel_index >= 5093) && (pixel_index <= 5132)) || ((pixel_index >= 5148) && (pixel_index <= 5177)) || ((pixel_index >= 5189) && (pixel_index <= 5230)) || ((pixel_index >= 5243) && (pixel_index <= 5273)) || ((pixel_index >= 5285) && (pixel_index <= 5328)) || ((pixel_index >= 5338) && (pixel_index <= 5369)) || ((pixel_index >= 5381) && (pixel_index <= 5465)) || ((pixel_index >= 5477) && (pixel_index <= 5561)) || ((pixel_index >= 5573) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 6041)) || (pixel_index >= 6053) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 23) begin
            if (((pixel_index >= 5) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 377)) || ((pixel_index >= 389) && (pixel_index <= 473)) || ((pixel_index >= 485) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 857)) || ((pixel_index >= 869) && (pixel_index <= 953)) || ((pixel_index >= 965) && (pixel_index <= 1049)) || ((pixel_index >= 1061) && (pixel_index <= 1145)) || ((pixel_index >= 1157) && (pixel_index <= 1241)) || ((pixel_index >= 1253) && (pixel_index <= 1337)) || ((pixel_index >= 1349) && (pixel_index <= 1433)) || ((pixel_index >= 1445) && (pixel_index <= 1529)) || ((pixel_index >= 1541) && (pixel_index <= 1625)) || ((pixel_index >= 1637) && (pixel_index <= 1721)) || ((pixel_index >= 1733) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2736)) || ((pixel_index >= 2738) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2832)) || ((pixel_index >= 2834) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2928)) || ((pixel_index >= 2938) && (pixel_index <= 2969)) || ((pixel_index >= 2981) && (pixel_index <= 3021)) || ((pixel_index >= 3035) && (pixel_index <= 3065)) || ((pixel_index >= 3077) && (pixel_index <= 3114)) || ((pixel_index >= 3132) && (pixel_index <= 3161)) || ((pixel_index >= 3173) && (pixel_index <= 3209)) || ((pixel_index >= 3229) && (pixel_index <= 3257)) || ((pixel_index >= 3269) && (pixel_index <= 3304)) || ((pixel_index >= 3325) && (pixel_index <= 3353)) || ((pixel_index >= 3365) && (pixel_index <= 3400)) || ((pixel_index >= 3422) && (pixel_index <= 3449)) || ((pixel_index >= 3461) && (pixel_index <= 3496)) || ((pixel_index >= 3518) && (pixel_index <= 3545)) || ((pixel_index >= 3557) && (pixel_index <= 3591)) || ((pixel_index >= 3614) && (pixel_index <= 3641)) || ((pixel_index >= 3653) && (pixel_index <= 3687)) || ((pixel_index >= 3710) && (pixel_index <= 3737)) || ((pixel_index >= 3749) && (pixel_index <= 3783)) || ((pixel_index >= 3806) && (pixel_index <= 3833)) || ((pixel_index >= 3845) && (pixel_index <= 3880)) || ((pixel_index >= 3902) && (pixel_index <= 3929)) || ((pixel_index >= 3941) && (pixel_index <= 3976)) || ((pixel_index >= 3998) && (pixel_index <= 4025)) || ((pixel_index >= 4037) && (pixel_index <= 4072)) || ((pixel_index >= 4094) && (pixel_index <= 4121)) || ((pixel_index >= 4133) && (pixel_index <= 4168)) || ((pixel_index >= 4190) && (pixel_index <= 4217)) || ((pixel_index >= 4229) && (pixel_index <= 4265)) || ((pixel_index >= 4285) && (pixel_index <= 4313)) || ((pixel_index >= 4325) && (pixel_index <= 4361)) || ((pixel_index >= 4381) && (pixel_index <= 4409)) || ((pixel_index >= 4421) && (pixel_index <= 4457)) || ((pixel_index >= 4477) && (pixel_index <= 4505)) || ((pixel_index >= 4517) && (pixel_index <= 4554)) || ((pixel_index >= 4572) && (pixel_index <= 4601)) || ((pixel_index >= 4613) && (pixel_index <= 4651)) || ((pixel_index >= 4668) && (pixel_index <= 4697)) || ((pixel_index >= 4709) && (pixel_index <= 4748)) || ((pixel_index >= 4763) && (pixel_index <= 4793)) || ((pixel_index >= 4805) && (pixel_index <= 4845)) || ((pixel_index >= 4857) && (pixel_index <= 4889)) || ((pixel_index >= 4901) && (pixel_index <= 4985)) || ((pixel_index >= 4997) && (pixel_index <= 5081)) || ((pixel_index >= 5093) && (pixel_index <= 5177)) || ((pixel_index >= 5189) && (pixel_index <= 5273)) || ((pixel_index >= 5285) && (pixel_index <= 5369)) || ((pixel_index >= 5381) && (pixel_index <= 5465)) || ((pixel_index >= 5477) && (pixel_index <= 5561)) || ((pixel_index >= 5573) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 6041)) || (pixel_index >= 6053) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 24) begin
            if (((pixel_index >= 5) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 377)) || ((pixel_index >= 389) && (pixel_index <= 473)) || ((pixel_index >= 485) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 857)) || ((pixel_index >= 869) && (pixel_index <= 953)) || ((pixel_index >= 965) && (pixel_index <= 1049)) || ((pixel_index >= 1061) && (pixel_index <= 1145)) || ((pixel_index >= 1157) && (pixel_index <= 1241)) || ((pixel_index >= 1253) && (pixel_index <= 1337)) || ((pixel_index >= 1349) && (pixel_index <= 1433)) || ((pixel_index >= 1445) && (pixel_index <= 1529)) || ((pixel_index >= 1541) && (pixel_index <= 1625)) || ((pixel_index >= 1637) && (pixel_index <= 1721)) || ((pixel_index >= 1733) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2060)) || ((pixel_index >= 2073) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2154)) || ((pixel_index >= 2170) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2248)) || ((pixel_index >= 2267) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2343)) || ((pixel_index >= 2363) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2439)) || ((pixel_index >= 2460) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2534)) || ((pixel_index >= 2556) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2630)) || ((pixel_index >= 2652) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2726)) || ((pixel_index >= 2749) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2822)) || ((pixel_index >= 2845) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2919)) || ((pixel_index >= 2942) && (pixel_index <= 2969)) || ((pixel_index >= 2981) && (pixel_index <= 3015)) || ((pixel_index >= 3038) && (pixel_index <= 3065)) || ((pixel_index >= 3077) && (pixel_index <= 3111)) || ((pixel_index >= 3134) && (pixel_index <= 3161)) || ((pixel_index >= 3173) && (pixel_index <= 3207)) || ((pixel_index >= 3230) && (pixel_index <= 3257)) || ((pixel_index >= 3269) && (pixel_index <= 3304)) || ((pixel_index >= 3326) && (pixel_index <= 3353)) || ((pixel_index >= 3365) && (pixel_index <= 3397)) || ((pixel_index >= 3421) && (pixel_index <= 3449)) || ((pixel_index >= 3461) && (pixel_index <= 3493)) || ((pixel_index >= 3495) && (pixel_index <= 3497)) || ((pixel_index >= 3517) && (pixel_index <= 3545)) || ((pixel_index >= 3557) && (pixel_index <= 3593)) || ((pixel_index >= 3612) && (pixel_index <= 3641)) || ((pixel_index >= 3653) && (pixel_index <= 3689)) || ((pixel_index >= 3707) && (pixel_index <= 3737)) || ((pixel_index >= 3749) && (pixel_index <= 3786)) || ((pixel_index >= 3802) && (pixel_index <= 3833)) || ((pixel_index >= 3845) && (pixel_index <= 3882)) || ((pixel_index >= 3897) && (pixel_index <= 3929)) || ((pixel_index >= 3941) && (pixel_index <= 3979)) || ((pixel_index >= 3991) && (pixel_index <= 4025)) || ((pixel_index >= 4037) && (pixel_index <= 4077)) || ((pixel_index >= 4085) && (pixel_index <= 4121)) || ((pixel_index >= 4133) && (pixel_index <= 4217)) || ((pixel_index >= 4229) && (pixel_index <= 4313)) || ((pixel_index >= 4325) && (pixel_index <= 4409)) || ((pixel_index >= 4421) && (pixel_index <= 4505)) || ((pixel_index >= 4517) && (pixel_index <= 4601)) || ((pixel_index >= 4613) && (pixel_index <= 4697)) || ((pixel_index >= 4709) && (pixel_index <= 4793)) || ((pixel_index >= 4805) && (pixel_index <= 4889)) || ((pixel_index >= 4901) && (pixel_index <= 4985)) || ((pixel_index >= 4997) && (pixel_index <= 5081)) || ((pixel_index >= 5093) && (pixel_index <= 5177)) || ((pixel_index >= 5189) && (pixel_index <= 5273)) || ((pixel_index >= 5285) && (pixel_index <= 5369)) || ((pixel_index >= 5381) && (pixel_index <= 5465)) || ((pixel_index >= 5477) && (pixel_index <= 5561)) || ((pixel_index >= 5573) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 6041)) || (pixel_index >= 6053) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 25) begin
            if (((pixel_index >= 5) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 377)) || ((pixel_index >= 389) && (pixel_index <= 473)) || ((pixel_index >= 485) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 857)) || ((pixel_index >= 869) && (pixel_index <= 953)) || ((pixel_index >= 965) && (pixel_index <= 1049)) || ((pixel_index >= 1061) && (pixel_index <= 1145)) || ((pixel_index >= 1157) && (pixel_index <= 1241)) || ((pixel_index >= 1253) && (pixel_index <= 1337)) || ((pixel_index >= 1349) && (pixel_index <= 1389)) || ((pixel_index >= 1396) && (pixel_index <= 1433)) || ((pixel_index >= 1445) && (pixel_index <= 1483)) || ((pixel_index >= 1494) && (pixel_index <= 1529)) || ((pixel_index >= 1541) && (pixel_index <= 1579)) || ((pixel_index >= 1591) && (pixel_index <= 1625)) || ((pixel_index >= 1637) && (pixel_index <= 1673)) || ((pixel_index >= 1689) && (pixel_index <= 1721)) || ((pixel_index >= 1733) && (pixel_index <= 1767)) || ((pixel_index >= 1786) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1862)) || ((pixel_index >= 1882) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 1958)) || ((pixel_index >= 1979) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2053)) || ((pixel_index >= 2076) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2149)) || ((pixel_index >= 2173) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2245)) || ((pixel_index >= 2269) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2341)) || ((pixel_index >= 2365) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2437)) || ((pixel_index >= 2461) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2533)) || ((pixel_index >= 2557) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2629)) || ((pixel_index >= 2653) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2726)) || ((pixel_index >= 2749) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2822)) || ((pixel_index >= 2845) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2918)) || ((pixel_index >= 2940) && (pixel_index <= 2969)) || ((pixel_index >= 2981) && (pixel_index <= 3014)) || ((pixel_index >= 3036) && (pixel_index <= 3065)) || ((pixel_index >= 3077) && (pixel_index <= 3111)) || ((pixel_index >= 3131) && (pixel_index <= 3161)) || ((pixel_index >= 3173) && (pixel_index <= 3207)) || ((pixel_index >= 3225) && (pixel_index <= 3257)) || ((pixel_index >= 3269) && (pixel_index <= 3304)) || ((pixel_index >= 3320) && (pixel_index <= 3353)) || ((pixel_index >= 3365) && (pixel_index <= 3401)) || ((pixel_index >= 3416) && (pixel_index <= 3449)) || ((pixel_index >= 3461) && (pixel_index <= 3497)) || ((pixel_index >= 3508) && (pixel_index <= 3510)) || ((pixel_index >= 3512) && (pixel_index <= 3545)) || ((pixel_index >= 3557) && (pixel_index <= 3595)) || ((pixel_index >= 3602) && (pixel_index <= 3607)) || ((pixel_index >= 3609) && (pixel_index <= 3641)) || ((pixel_index >= 3653) && (pixel_index <= 3703)) || ((pixel_index >= 3705) && (pixel_index <= 3737)) || ((pixel_index >= 3749) && (pixel_index <= 3833)) || ((pixel_index >= 3845) && (pixel_index <= 3929)) || ((pixel_index >= 3941) && (pixel_index <= 4025)) || ((pixel_index >= 4037) && (pixel_index <= 4121)) || ((pixel_index >= 4133) && (pixel_index <= 4217)) || ((pixel_index >= 4229) && (pixel_index <= 4313)) || ((pixel_index >= 4325) && (pixel_index <= 4409)) || ((pixel_index >= 4421) && (pixel_index <= 4505)) || ((pixel_index >= 4517) && (pixel_index <= 4601)) || ((pixel_index >= 4613) && (pixel_index <= 4697)) || ((pixel_index >= 4709) && (pixel_index <= 4793)) || ((pixel_index >= 4805) && (pixel_index <= 4889)) || ((pixel_index >= 4901) && (pixel_index <= 4985)) || ((pixel_index >= 4997) && (pixel_index <= 5081)) || ((pixel_index >= 5093) && (pixel_index <= 5177)) || ((pixel_index >= 5189) && (pixel_index <= 5273)) || ((pixel_index >= 5285) && (pixel_index <= 5369)) || ((pixel_index >= 5381) && (pixel_index <= 5465)) || ((pixel_index >= 5477) && (pixel_index <= 5561)) || ((pixel_index >= 5573) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 6041)) || (pixel_index >= 6053) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 26) begin
            if (((pixel_index >= 5) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 377)) || ((pixel_index >= 389) && (pixel_index <= 473)) || ((pixel_index >= 485) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 857)) || ((pixel_index >= 869) && (pixel_index <= 953)) || ((pixel_index >= 965) && (pixel_index <= 1049)) || ((pixel_index >= 1061) && (pixel_index <= 1145)) || ((pixel_index >= 1157) && (pixel_index <= 1241)) || ((pixel_index >= 1253) && (pixel_index <= 1337)) || ((pixel_index >= 1349) && (pixel_index <= 1433)) || ((pixel_index >= 1445) && (pixel_index <= 1486)) || ((pixel_index >= 1493) && (pixel_index <= 1529)) || ((pixel_index >= 1541) && (pixel_index <= 1580)) || ((pixel_index >= 1591) && (pixel_index <= 1625)) || ((pixel_index >= 1637) && (pixel_index <= 1675)) || ((pixel_index >= 1688) && (pixel_index <= 1721)) || ((pixel_index >= 1733) && (pixel_index <= 1770)) || ((pixel_index >= 1785) && (pixel_index <= 1787)) || ((pixel_index >= 1790) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1865)) || pixel_index == 1882 || ((pixel_index >= 1885) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 1960)) || ((pixel_index >= 1980) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2055)) || ((pixel_index >= 2075) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2151)) || ((pixel_index >= 2172) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2246)) || ((pixel_index >= 2269) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2342)) || ((pixel_index >= 2366) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2438)) || ((pixel_index >= 2462) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2533)) || ((pixel_index >= 2558) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2629)) || ((pixel_index >= 2655) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2725)) || ((pixel_index >= 2751) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2821)) || ((pixel_index >= 2847) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2917)) || ((pixel_index >= 2943) && (pixel_index <= 2969)) || ((pixel_index >= 2981) && (pixel_index <= 3014)) || ((pixel_index >= 3039) && (pixel_index <= 3065)) || ((pixel_index >= 3077) && (pixel_index <= 3110)) || ((pixel_index >= 3134) && (pixel_index <= 3161)) || ((pixel_index >= 3173) && (pixel_index <= 3207)) || ((pixel_index >= 3229) && (pixel_index <= 3257)) || ((pixel_index >= 3269) && (pixel_index <= 3304)) || ((pixel_index >= 3324) && (pixel_index <= 3353)) || ((pixel_index >= 3365) && (pixel_index <= 3401)) || ((pixel_index >= 3419) && (pixel_index <= 3449)) || ((pixel_index >= 3461) && (pixel_index <= 3497)) || ((pixel_index >= 3514) && (pixel_index <= 3545)) || ((pixel_index >= 3557) && (pixel_index <= 3594)) || ((pixel_index >= 3608) && (pixel_index <= 3641)) || ((pixel_index >= 3653) && (pixel_index <= 3691)) || ((pixel_index >= 3702) && (pixel_index <= 3737)) || ((pixel_index >= 3749) && (pixel_index <= 3791)) || ((pixel_index >= 3793) && (pixel_index <= 3833)) || ((pixel_index >= 3845) && (pixel_index <= 3929)) || ((pixel_index >= 3941) && (pixel_index <= 4025)) || ((pixel_index >= 4037) && (pixel_index <= 4121)) || ((pixel_index >= 4133) && (pixel_index <= 4217)) || ((pixel_index >= 4229) && (pixel_index <= 4313)) || ((pixel_index >= 4325) && (pixel_index <= 4409)) || ((pixel_index >= 4421) && (pixel_index <= 4505)) || ((pixel_index >= 4517) && (pixel_index <= 4601)) || ((pixel_index >= 4613) && (pixel_index <= 4697)) || ((pixel_index >= 4709) && (pixel_index <= 4793)) || ((pixel_index >= 4805) && (pixel_index <= 4889)) || ((pixel_index >= 4901) && (pixel_index <= 4985)) || ((pixel_index >= 4997) && (pixel_index <= 5081)) || ((pixel_index >= 5093) && (pixel_index <= 5177)) || ((pixel_index >= 5189) && (pixel_index <= 5273)) || ((pixel_index >= 5285) && (pixel_index <= 5369)) || ((pixel_index >= 5381) && (pixel_index <= 5465)) || ((pixel_index >= 5477) && (pixel_index <= 5561)) || ((pixel_index >= 5573) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 6041)) || (pixel_index >= 6053) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 27) begin
            if (((pixel_index >= 5) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 377)) || ((pixel_index >= 389) && (pixel_index <= 473)) || ((pixel_index >= 485) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 857)) || ((pixel_index >= 869) && (pixel_index <= 953)) || ((pixel_index >= 965) && (pixel_index <= 1049)) || ((pixel_index >= 1061) && (pixel_index <= 1145)) || ((pixel_index >= 1157) && (pixel_index <= 1241)) || ((pixel_index >= 1253) && (pixel_index <= 1337)) || ((pixel_index >= 1349) && (pixel_index <= 1433)) || ((pixel_index >= 1445) && (pixel_index <= 1529)) || ((pixel_index >= 1541) && (pixel_index <= 1625)) || ((pixel_index >= 1637) && (pixel_index <= 1721)) || ((pixel_index >= 1733) && (pixel_index <= 1777)) || ((pixel_index >= 1786) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1871)) || ((pixel_index >= 1883) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 1963)) || ((pixel_index >= 1965) && (pixel_index <= 1966)) || ((pixel_index >= 1980) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2059)) || ((pixel_index >= 2077) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2155)) || ((pixel_index >= 2174) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2250)) || ((pixel_index >= 2270) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2346)) || ((pixel_index >= 2367) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2441)) || ((pixel_index >= 2463) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2536)) || ((pixel_index >= 2560) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2632)) || ((pixel_index >= 2656) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2727)) || ((pixel_index >= 2753) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2823)) || ((pixel_index >= 2849) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2919)) || ((pixel_index >= 2945) && (pixel_index <= 2969)) || ((pixel_index >= 2981) && (pixel_index <= 3015)) || ((pixel_index >= 3041) && (pixel_index <= 3065)) || ((pixel_index >= 3077) && (pixel_index <= 3111)) || ((pixel_index >= 3137) && (pixel_index <= 3161)) || ((pixel_index >= 3173) && (pixel_index <= 3207)) || ((pixel_index >= 3233) && (pixel_index <= 3257)) || ((pixel_index >= 3269) && (pixel_index <= 3303)) || ((pixel_index >= 3329) && (pixel_index <= 3353)) || ((pixel_index >= 3365) && (pixel_index <= 3400)) || ((pixel_index >= 3425) && (pixel_index <= 3449)) || ((pixel_index >= 3461) && (pixel_index <= 3497)) || ((pixel_index >= 3520) && (pixel_index <= 3545)) || ((pixel_index >= 3557) && (pixel_index <= 3594)) || ((pixel_index >= 3614) && (pixel_index <= 3641)) || ((pixel_index >= 3653) && (pixel_index <= 3690)) || ((pixel_index >= 3709) && (pixel_index <= 3737)) || ((pixel_index >= 3749) && (pixel_index <= 3788)) || ((pixel_index >= 3805) && (pixel_index <= 3833)) || ((pixel_index >= 3845) && (pixel_index <= 3885)) || ((pixel_index >= 3900) && (pixel_index <= 3929)) || ((pixel_index >= 3941) && (pixel_index <= 3983)) || ((pixel_index >= 3995) && (pixel_index <= 4025)) || ((pixel_index >= 4037) && (pixel_index <= 4081)) || ((pixel_index >= 4089) && (pixel_index <= 4121)) || ((pixel_index >= 4133) && (pixel_index <= 4217)) || ((pixel_index >= 4229) && (pixel_index <= 4313)) || ((pixel_index >= 4325) && (pixel_index <= 4409)) || ((pixel_index >= 4421) && (pixel_index <= 4505)) || ((pixel_index >= 4517) && (pixel_index <= 4601)) || ((pixel_index >= 4613) && (pixel_index <= 4697)) || ((pixel_index >= 4709) && (pixel_index <= 4793)) || ((pixel_index >= 4805) && (pixel_index <= 4889)) || ((pixel_index >= 4901) && (pixel_index <= 4985)) || ((pixel_index >= 4997) && (pixel_index <= 5081)) || ((pixel_index >= 5093) && (pixel_index <= 5177)) || ((pixel_index >= 5189) && (pixel_index <= 5273)) || ((pixel_index >= 5285) && (pixel_index <= 5369)) || ((pixel_index >= 5381) && (pixel_index <= 5465)) || ((pixel_index >= 5477) && (pixel_index <= 5561)) || ((pixel_index >= 5573) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 6041)) || (pixel_index >= 6053) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 28) begin
            if (((pixel_index >= 5) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 377)) || ((pixel_index >= 389) && (pixel_index <= 473)) || ((pixel_index >= 485) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 857)) || ((pixel_index >= 869) && (pixel_index <= 953)) || ((pixel_index >= 965) && (pixel_index <= 1049)) || ((pixel_index >= 1061) && (pixel_index <= 1145)) || ((pixel_index >= 1157) && (pixel_index <= 1241)) || ((pixel_index >= 1253) && (pixel_index <= 1337)) || ((pixel_index >= 1349) && (pixel_index <= 1433)) || ((pixel_index >= 1445) && (pixel_index <= 1529)) || ((pixel_index >= 1541) && (pixel_index <= 1625)) || ((pixel_index >= 1637) && (pixel_index <= 1721)) || ((pixel_index >= 1733) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2068)) || ((pixel_index >= 2075) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2161)) || ((pixel_index >= 2173) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2255)) || ((pixel_index >= 2270) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2349)) || ((pixel_index >= 2367) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2444)) || ((pixel_index >= 2463) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2539)) || ((pixel_index >= 2561) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2634)) || ((pixel_index >= 2658) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2729)) || ((pixel_index >= 2754) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2825)) || ((pixel_index >= 2851) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2921)) || ((pixel_index >= 2947) && (pixel_index <= 2969)) || ((pixel_index >= 2981) && (pixel_index <= 3016)) || ((pixel_index >= 3043) && (pixel_index <= 3065)) || ((pixel_index >= 3077) && (pixel_index <= 3112)) || ((pixel_index >= 3139) && (pixel_index <= 3161)) || ((pixel_index >= 3173) && (pixel_index <= 3208)) || ((pixel_index >= 3235) && (pixel_index <= 3257)) || ((pixel_index >= 3269) && (pixel_index <= 3304)) || ((pixel_index >= 3331) && (pixel_index <= 3353)) || ((pixel_index >= 3365) && (pixel_index <= 3400)) || ((pixel_index >= 3427) && (pixel_index <= 3449)) || ((pixel_index >= 3461) && (pixel_index <= 3497)) || ((pixel_index >= 3522) && (pixel_index <= 3545)) || ((pixel_index >= 3557) && (pixel_index <= 3593)) || ((pixel_index >= 3618) && (pixel_index <= 3641)) || ((pixel_index >= 3653) && (pixel_index <= 3689)) || ((pixel_index >= 3713) && (pixel_index <= 3737)) || ((pixel_index >= 3749) && (pixel_index <= 3785)) || ((pixel_index >= 3809) && (pixel_index <= 3833)) || ((pixel_index >= 3845) && (pixel_index <= 3882)) || ((pixel_index >= 3904) && (pixel_index <= 3929)) || ((pixel_index >= 3941) && (pixel_index <= 3979)) || ((pixel_index >= 4000) && (pixel_index <= 4025)) || ((pixel_index >= 4037) && (pixel_index <= 4076)) || ((pixel_index >= 4095) && (pixel_index <= 4121)) || ((pixel_index >= 4133) && (pixel_index <= 4173)) || ((pixel_index >= 4190) && (pixel_index <= 4217)) || ((pixel_index >= 4229) && (pixel_index <= 4271)) || ((pixel_index >= 4285) && (pixel_index <= 4313)) || ((pixel_index >= 4325) && (pixel_index <= 4368)) || ((pixel_index >= 4379) && (pixel_index <= 4409)) || ((pixel_index >= 4421) && (pixel_index <= 4465)) || ((pixel_index >= 4473) && (pixel_index <= 4505)) || ((pixel_index >= 4517) && (pixel_index <= 4601)) || ((pixel_index >= 4613) && (pixel_index <= 4697)) || ((pixel_index >= 4709) && (pixel_index <= 4793)) || ((pixel_index >= 4805) && (pixel_index <= 4889)) || ((pixel_index >= 4901) && (pixel_index <= 4985)) || ((pixel_index >= 4997) && (pixel_index <= 5081)) || ((pixel_index >= 5093) && (pixel_index <= 5177)) || ((pixel_index >= 5189) && (pixel_index <= 5273)) || ((pixel_index >= 5285) && (pixel_index <= 5369)) || ((pixel_index >= 5381) && (pixel_index <= 5465)) || ((pixel_index >= 5477) && (pixel_index <= 5561)) || ((pixel_index >= 5573) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 6041)) || (pixel_index >= 6053) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 29) begin
            if (((pixel_index >= 5) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 377)) || ((pixel_index >= 389) && (pixel_index <= 473)) || ((pixel_index >= 485) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 857)) || ((pixel_index >= 869) && (pixel_index <= 953)) || ((pixel_index >= 965) && (pixel_index <= 1049)) || ((pixel_index >= 1061) && (pixel_index <= 1145)) || ((pixel_index >= 1157) && (pixel_index <= 1241)) || ((pixel_index >= 1253) && (pixel_index <= 1337)) || ((pixel_index >= 1349) && (pixel_index <= 1433)) || ((pixel_index >= 1445) && (pixel_index <= 1529)) || ((pixel_index >= 1541) && (pixel_index <= 1625)) || ((pixel_index >= 1637) && (pixel_index <= 1721)) || ((pixel_index >= 1733) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2163)) || ((pixel_index >= 2166) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2255)) || ((pixel_index >= 2265) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2349)) || ((pixel_index >= 2363) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2444)) || ((pixel_index >= 2461) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2539)) || ((pixel_index >= 2558) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2635)) || ((pixel_index >= 2655) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2730)) || ((pixel_index >= 2752) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2825)) || ((pixel_index >= 2849) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2920)) || ((pixel_index >= 2946) && (pixel_index <= 2969)) || ((pixel_index >= 2981) && (pixel_index <= 3016)) || ((pixel_index >= 3042) && (pixel_index <= 3065)) || ((pixel_index >= 3077) && (pixel_index <= 3112)) || ((pixel_index >= 3138) && (pixel_index <= 3161)) || ((pixel_index >= 3173) && (pixel_index <= 3208)) || ((pixel_index >= 3235) && (pixel_index <= 3257)) || ((pixel_index >= 3269) && (pixel_index <= 3304)) || ((pixel_index >= 3331) && (pixel_index <= 3353)) || ((pixel_index >= 3365) && (pixel_index <= 3400)) || ((pixel_index >= 3427) && (pixel_index <= 3449)) || ((pixel_index >= 3461) && (pixel_index <= 3496)) || ((pixel_index >= 3523) && (pixel_index <= 3545)) || ((pixel_index >= 3557) && (pixel_index <= 3593)) || ((pixel_index >= 3618) && (pixel_index <= 3641)) || ((pixel_index >= 3653) && (pixel_index <= 3689)) || ((pixel_index >= 3714) && (pixel_index <= 3737)) || ((pixel_index >= 3749) && (pixel_index <= 3785)) || ((pixel_index >= 3809) && (pixel_index <= 3833)) || ((pixel_index >= 3845) && (pixel_index <= 3882)) || ((pixel_index >= 3904) && (pixel_index <= 3929)) || ((pixel_index >= 3941) && (pixel_index <= 3978)) || ((pixel_index >= 3999) && (pixel_index <= 4025)) || ((pixel_index >= 4037) && (pixel_index <= 4075)) || ((pixel_index >= 4094) && (pixel_index <= 4121)) || ((pixel_index >= 4133) && (pixel_index <= 4172)) || ((pixel_index >= 4189) && (pixel_index <= 4217)) || ((pixel_index >= 4229) && (pixel_index <= 4268)) || ((pixel_index >= 4283) && (pixel_index <= 4284)) || ((pixel_index >= 4286) && (pixel_index <= 4313)) || ((pixel_index >= 4325) && (pixel_index <= 4365)) || ((pixel_index >= 4378) && (pixel_index <= 4381)) || ((pixel_index >= 4383) && (pixel_index <= 4409)) || ((pixel_index >= 4421) && (pixel_index <= 4462)) || ((pixel_index >= 4473) && (pixel_index <= 4478)) || ((pixel_index >= 4480) && (pixel_index <= 4505)) || ((pixel_index >= 4517) && (pixel_index <= 4560)) || ((pixel_index >= 4567) && (pixel_index <= 4601)) || ((pixel_index >= 4613) && (pixel_index <= 4697)) || ((pixel_index >= 4709) && (pixel_index <= 4793)) || ((pixel_index >= 4805) && (pixel_index <= 4889)) || ((pixel_index >= 4901) && (pixel_index <= 4985)) || ((pixel_index >= 4997) && (pixel_index <= 5081)) || ((pixel_index >= 5093) && (pixel_index <= 5177)) || ((pixel_index >= 5189) && (pixel_index <= 5273)) || ((pixel_index >= 5285) && (pixel_index <= 5369)) || ((pixel_index >= 5381) && (pixel_index <= 5465)) || ((pixel_index >= 5477) && (pixel_index <= 5561)) || ((pixel_index >= 5573) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 6041)) || (pixel_index >= 6053) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 30) begin
            if (((pixel_index >= 5) && (pixel_index <= 28)) || ((pixel_index >= 101) && (pixel_index <= 129)) || ((pixel_index >= 197) && (pixel_index <= 233)) || ((pixel_index >= 293) && (pixel_index <= 337)) || ((pixel_index >= 343) && (pixel_index <= 348)) || ((pixel_index >= 389) && (pixel_index <= 465)) || pixel_index == 473 || ((pixel_index >= 485) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 857)) || ((pixel_index >= 869) && (pixel_index <= 953)) || ((pixel_index >= 965) && (pixel_index <= 1049)) || ((pixel_index >= 1061) && (pixel_index <= 1145)) || ((pixel_index >= 1157) && (pixel_index <= 1241)) || ((pixel_index >= 1253) && (pixel_index <= 1337)) || ((pixel_index >= 1349) && (pixel_index <= 1433)) || ((pixel_index >= 1445) && (pixel_index <= 1529)) || ((pixel_index >= 1541) && (pixel_index <= 1625)) || ((pixel_index >= 1637) && (pixel_index <= 1721)) || ((pixel_index >= 1733) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2260)) || ((pixel_index >= 2262) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2349)) || ((pixel_index >= 2361) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2443)) || ((pixel_index >= 2458) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2538)) || ((pixel_index >= 2556) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2633)) || ((pixel_index >= 2653) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2728)) || ((pixel_index >= 2751) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2824)) || ((pixel_index >= 2847) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2919)) || ((pixel_index >= 2944) && (pixel_index <= 2969)) || ((pixel_index >= 2981) && (pixel_index <= 3015)) || ((pixel_index >= 3040) && (pixel_index <= 3065)) || ((pixel_index >= 3077) && (pixel_index <= 3111)) || ((pixel_index >= 3136) && (pixel_index <= 3161)) || ((pixel_index >= 3173) && (pixel_index <= 3207)) || ((pixel_index >= 3233) && (pixel_index <= 3257)) || ((pixel_index >= 3269) && (pixel_index <= 3303)) || ((pixel_index >= 3329) && (pixel_index <= 3353)) || ((pixel_index >= 3365) && (pixel_index <= 3399)) || ((pixel_index >= 3425) && (pixel_index <= 3449)) || ((pixel_index >= 3461) && (pixel_index <= 3495)) || ((pixel_index >= 3520) && (pixel_index <= 3545)) || ((pixel_index >= 3557) && (pixel_index <= 3591)) || ((pixel_index >= 3616) && (pixel_index <= 3641)) || ((pixel_index >= 3653) && (pixel_index <= 3687)) || ((pixel_index >= 3712) && (pixel_index <= 3737)) || ((pixel_index >= 3749) && (pixel_index <= 3783)) || ((pixel_index >= 3807) && (pixel_index <= 3833)) || ((pixel_index >= 3845) && (pixel_index <= 3880)) || ((pixel_index >= 3903) && (pixel_index <= 3929)) || ((pixel_index >= 3941) && (pixel_index <= 3976)) || ((pixel_index >= 3998) && (pixel_index <= 4025)) || ((pixel_index >= 4037) && (pixel_index <= 4073)) || ((pixel_index >= 4093) && (pixel_index <= 4121)) || ((pixel_index >= 4133) && (pixel_index <= 4169)) || ((pixel_index >= 4189) && (pixel_index <= 4217)) || ((pixel_index >= 4229) && (pixel_index <= 4266)) || ((pixel_index >= 4284) && (pixel_index <= 4313)) || ((pixel_index >= 4325) && (pixel_index <= 4363)) || ((pixel_index >= 4378) && (pixel_index <= 4409)) || ((pixel_index >= 4421) && (pixel_index <= 4461)) || ((pixel_index >= 4473) && (pixel_index <= 4505)) || ((pixel_index >= 4517) && (pixel_index <= 4558)) || ((pixel_index >= 4567) && (pixel_index <= 4601)) || ((pixel_index >= 4613) && (pixel_index <= 4697)) || ((pixel_index >= 4709) && (pixel_index <= 4793)) || ((pixel_index >= 4805) && (pixel_index <= 4889)) || ((pixel_index >= 4901) && (pixel_index <= 4985)) || ((pixel_index >= 4997) && (pixel_index <= 5081)) || ((pixel_index >= 5093) && (pixel_index <= 5177)) || ((pixel_index >= 5189) && (pixel_index <= 5273)) || ((pixel_index >= 5285) && (pixel_index <= 5369)) || ((pixel_index >= 5381) && (pixel_index <= 5465)) || ((pixel_index >= 5477) && (pixel_index <= 5561)) || ((pixel_index >= 5573) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 6041)) || (pixel_index >= 6053) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 31) begin
            oled_data = 0;
            done = 1;
        end
    end
    
endmodule

module o_win_anim(input frame_rate, input start, input [12:0] pixel_index, output reg done, output reg [15:0] oled_data);
    reg [15:0] frame_count = 0;
    
    always @ (posedge frame_rate) begin
        if (start) frame_count <= (frame_count == 31) ? 31 : frame_count + 1;
        else frame_count <= 0;
    end
   
    // animation for O win (1v1 mode) or player lose (AI mode)
    // Remilia dropping teacup
    always @ (*) begin
        if (frame_count <= 30) done = 0;
        if (frame_count == 0) oled_data = 0;
        else if (frame_count == 1) begin
            if (((pixel_index >= 5) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 377)) || ((pixel_index >= 389) && (pixel_index <= 473)) || ((pixel_index >= 485) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 809)) || ((pixel_index >= 820) && (pixel_index <= 827)) || ((pixel_index >= 829) && (pixel_index <= 857)) || ((pixel_index >= 869) && (pixel_index <= 903)) || ((pixel_index >= 918) && (pixel_index <= 922)) || ((pixel_index >= 925) && (pixel_index <= 953)) || ((pixel_index >= 965) && (pixel_index <= 998)) || ((pixel_index >= 1015) && (pixel_index <= 1017)) || ((pixel_index >= 1021) && (pixel_index <= 1049)) || ((pixel_index >= 1061) && (pixel_index <= 1094)) || ((pixel_index >= 1118) && (pixel_index <= 1145)) || ((pixel_index >= 1157) && (pixel_index <= 1189)) || ((pixel_index >= 1214) && (pixel_index <= 1241)) || ((pixel_index >= 1253) && (pixel_index <= 1285)) || ((pixel_index >= 1311) && (pixel_index <= 1337)) || ((pixel_index >= 1349) && (pixel_index <= 1381)) || ((pixel_index >= 1407) && (pixel_index <= 1433)) || ((pixel_index >= 1445) && (pixel_index <= 1477)) || ((pixel_index >= 1504) && (pixel_index <= 1529)) || ((pixel_index >= 1541) && (pixel_index <= 1573)) || ((pixel_index >= 1597) && (pixel_index <= 1625)) || ((pixel_index >= 1637) && (pixel_index <= 1669)) || ((pixel_index >= 1693) && (pixel_index <= 1721)) || ((pixel_index >= 1733) && (pixel_index <= 1763)) || ((pixel_index >= 1789) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1858)) || ((pixel_index >= 1884) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 1953)) || ((pixel_index >= 1978) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2050)) || ((pixel_index >= 2075) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2147)) || ((pixel_index >= 2171) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2245)) || ((pixel_index >= 2265) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2342)) || ((pixel_index >= 2360) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2437)) || ((pixel_index >= 2456) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2532)) || ((pixel_index >= 2552) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2629)) || ((pixel_index >= 2649) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2727)) || ((pixel_index >= 2744) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2824)) || ((pixel_index >= 2838) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2923)) || ((pixel_index >= 2930) && (pixel_index <= 2969)) || ((pixel_index >= 2981) && (pixel_index <= 3019)) || ((pixel_index >= 3026) && (pixel_index <= 3065)) || ((pixel_index >= 3077) && (pixel_index <= 3084)) || ((pixel_index >= 3087) && (pixel_index <= 3110)) || ((pixel_index >= 3125) && (pixel_index <= 3161)) || ((pixel_index >= 3173) && (pixel_index <= 3179)) || ((pixel_index >= 3185) && (pixel_index <= 3204)) || ((pixel_index >= 3224) && (pixel_index <= 3257)) || ((pixel_index >= 3269) && (pixel_index <= 3274)) || ((pixel_index >= 3283) && (pixel_index <= 3299)) || ((pixel_index >= 3321) && (pixel_index <= 3340)) || ((pixel_index >= 3342) && (pixel_index <= 3353)) || ((pixel_index >= 3365) && (pixel_index <= 3369)) || ((pixel_index >= 3381) && (pixel_index <= 3395)) || ((pixel_index >= 3418) && (pixel_index <= 3435)) || ((pixel_index >= 3439) && (pixel_index <= 3449)) || ((pixel_index >= 3461) && (pixel_index <= 3465)) || ((pixel_index >= 3478) && (pixel_index <= 3490)) || ((pixel_index >= 3515) && (pixel_index <= 3529)) || ((pixel_index >= 3536) && (pixel_index <= 3545)) || ((pixel_index >= 3557) && (pixel_index <= 3560)) || ((pixel_index >= 3576) && (pixel_index <= 3586)) || ((pixel_index >= 3611) && (pixel_index <= 3623)) || ((pixel_index >= 3633) && (pixel_index <= 3641)) || ((pixel_index >= 3653) && (pixel_index <= 3655)) || ((pixel_index >= 3674) && (pixel_index <= 3682)) || ((pixel_index >= 3708) && (pixel_index <= 3717)) || ((pixel_index >= 3729) && (pixel_index <= 3737)) || ((pixel_index >= 3749) && (pixel_index <= 3750)) || ((pixel_index >= 3804) && (pixel_index <= 3811)) || ((pixel_index >= 3826) && (pixel_index <= 3833)) || ((pixel_index >= 3902) && (pixel_index <= 3905)) || ((pixel_index >= 3923) && (pixel_index <= 3929)) || ((pixel_index >= 4020) && (pixel_index <= 4025)) || ((pixel_index >= 4066) && (pixel_index <= 4067)) || ((pixel_index >= 4117) && (pixel_index <= 4121)) || pixel_index == 4139 || pixel_index == 4143 || ((pixel_index >= 4161) && (pixel_index <= 4163)) || ((pixel_index >= 4214) && (pixel_index <= 4217)) || ((pixel_index >= 4234) && (pixel_index <= 4236)) || ((pixel_index >= 4238) && (pixel_index <= 4241)) || ((pixel_index >= 4255) && (pixel_index <= 4259)) || ((pixel_index >= 4312) && (pixel_index <= 4313)) || ((pixel_index >= 4330) && (pixel_index <= 4338)) || ((pixel_index >= 4341) && (pixel_index <= 4345)) || ((pixel_index >= 4350) && (pixel_index <= 4356)) || pixel_index == 4379 || pixel_index == 4409 || ((pixel_index >= 4425) && (pixel_index <= 4442)) || ((pixel_index >= 4444) && (pixel_index <= 4452)) || ((pixel_index >= 4475) && (pixel_index <= 4476)) || pixel_index == 4483 || ((pixel_index >= 4490) && (pixel_index <= 4492)) || pixel_index == 4495 || ((pixel_index >= 4517) && (pixel_index <= 4548)) || ((pixel_index >= 4571) && (pixel_index <= 4573)) || ((pixel_index >= 4577) && (pixel_index <= 4581)) || ((pixel_index >= 4584) && (pixel_index <= 4588)) || ((pixel_index >= 4590) && (pixel_index <= 4592)) || ((pixel_index >= 4613) && (pixel_index <= 4644)) || ((pixel_index >= 4667) && (pixel_index <= 4689)) || ((pixel_index >= 4709) && (pixel_index <= 4740)) || ((pixel_index >= 4763) && (pixel_index <= 4786)) || pixel_index == 4792 || ((pixel_index >= 4805) && (pixel_index <= 4836)) || ((pixel_index >= 4859) && (pixel_index <= 4882)) || ((pixel_index >= 4885) && (pixel_index <= 4889)) || ((pixel_index >= 4901) && (pixel_index <= 4933)) || ((pixel_index >= 4949) && (pixel_index <= 4950)) || ((pixel_index >= 4955) && (pixel_index <= 4985)) || ((pixel_index >= 4997) && (pixel_index <= 5029)) || ((pixel_index >= 5045) && (pixel_index <= 5046)) || ((pixel_index >= 5050) && (pixel_index <= 5081)) || ((pixel_index >= 5093) && (pixel_index <= 5125)) || ((pixel_index >= 5141) && (pixel_index <= 5177)) || ((pixel_index >= 5189) && (pixel_index <= 5221)) || ((pixel_index >= 5237) && (pixel_index <= 5273)) || ((pixel_index >= 5285) && (pixel_index <= 5316)) || ((pixel_index >= 5333) && (pixel_index <= 5369)) || ((pixel_index >= 5381) && (pixel_index <= 5411)) || ((pixel_index >= 5430) && (pixel_index <= 5465)) || ((pixel_index >= 5477) && (pixel_index <= 5508)) || ((pixel_index >= 5526) && (pixel_index <= 5561)) || ((pixel_index >= 5573) && (pixel_index <= 5603)) || ((pixel_index >= 5622) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5700)) || ((pixel_index >= 5718) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5795)) || ((pixel_index >= 5814) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5891)) || ((pixel_index >= 5910) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 5986)) || ((pixel_index >= 6007) && (pixel_index <= 6041)) || ((pixel_index >= 6053) && (pixel_index <= 6082)) || (pixel_index >= 6103) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 2) begin
            if (((pixel_index >= 5) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 377)) || ((pixel_index >= 389) && (pixel_index <= 473)) || ((pixel_index >= 485) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 857)) || ((pixel_index >= 869) && (pixel_index <= 904)) || ((pixel_index >= 917) && (pixel_index <= 953)) || ((pixel_index >= 965) && (pixel_index <= 999)) || ((pixel_index >= 1014) && (pixel_index <= 1049)) || ((pixel_index >= 1061) && (pixel_index <= 1094)) || ((pixel_index >= 1111) && (pixel_index <= 1114)) || ((pixel_index >= 1117) && (pixel_index <= 1145)) || ((pixel_index >= 1157) && (pixel_index <= 1189)) || pixel_index == 1208 || ((pixel_index >= 1213) && (pixel_index <= 1241)) || ((pixel_index >= 1253) && (pixel_index <= 1285)) || ((pixel_index >= 1309) && (pixel_index <= 1337)) || ((pixel_index >= 1349) && (pixel_index <= 1381)) || ((pixel_index >= 1405) && (pixel_index <= 1433)) || ((pixel_index >= 1445) && (pixel_index <= 1477)) || ((pixel_index >= 1502) && (pixel_index <= 1529)) || ((pixel_index >= 1541) && (pixel_index <= 1573)) || ((pixel_index >= 1598) && (pixel_index <= 1625)) || ((pixel_index >= 1637) && (pixel_index <= 1669)) || ((pixel_index >= 1695) && (pixel_index <= 1721)) || ((pixel_index >= 1733) && (pixel_index <= 1764)) || ((pixel_index >= 1791) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1859)) || ((pixel_index >= 1884) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 1954)) || ((pixel_index >= 1980) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2049)) || pixel_index == 2073 || ((pixel_index >= 2076) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2146)) || ((pixel_index >= 2170) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2245)) || ((pixel_index >= 2266) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2341)) || ((pixel_index >= 2360) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2437)) || ((pixel_index >= 2456) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2532)) || ((pixel_index >= 2551) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2628)) || ((pixel_index >= 2648) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2725)) || ((pixel_index >= 2744) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2823)) || ((pixel_index >= 2839) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2920)) || ((pixel_index >= 2933) && (pixel_index <= 2969)) || ((pixel_index >= 2981) && (pixel_index <= 2986)) || ((pixel_index >= 2988) && (pixel_index <= 3018)) || ((pixel_index >= 3025) && (pixel_index <= 3065)) || ((pixel_index >= 3077) && (pixel_index <= 3081)) || ((pixel_index >= 3085) && (pixel_index <= 3113)) || ((pixel_index >= 3122) && (pixel_index <= 3161)) || ((pixel_index >= 3173) && (pixel_index <= 3177)) || ((pixel_index >= 3182) && (pixel_index <= 3204)) || ((pixel_index >= 3220) && (pixel_index <= 3257)) || ((pixel_index >= 3269) && (pixel_index <= 3272)) || ((pixel_index >= 3280) && (pixel_index <= 3299)) || ((pixel_index >= 3319) && (pixel_index <= 3353)) || ((pixel_index >= 3365) && (pixel_index <= 3367)) || ((pixel_index >= 3378) && (pixel_index <= 3395)) || ((pixel_index >= 3416) && (pixel_index <= 3434)) || ((pixel_index >= 3436) && (pixel_index <= 3449)) || ((pixel_index >= 3461) && (pixel_index <= 3462)) || ((pixel_index >= 3475) && (pixel_index <= 3490)) || ((pixel_index >= 3513) && (pixel_index <= 3529)) || ((pixel_index >= 3532) && (pixel_index <= 3545)) || pixel_index == 3557 || ((pixel_index >= 3573) && (pixel_index <= 3586)) || ((pixel_index >= 3610) && (pixel_index <= 3622)) || ((pixel_index >= 3629) && (pixel_index <= 3641)) || ((pixel_index >= 3670) && (pixel_index <= 3681)) || ((pixel_index >= 3706) && (pixel_index <= 3716)) || ((pixel_index >= 3726) && (pixel_index <= 3737)) || ((pixel_index >= 3769) && (pixel_index <= 3771)) || ((pixel_index >= 3775) && (pixel_index <= 3777)) || ((pixel_index >= 3803) && (pixel_index <= 3810)) || ((pixel_index >= 3822) && (pixel_index <= 3833)) || ((pixel_index >= 3899) && (pixel_index <= 3905)) || ((pixel_index >= 3919) && (pixel_index <= 3929)) || ((pixel_index >= 4016) && (pixel_index <= 4025)) || pixel_index == 4066 || ((pixel_index >= 4112) && (pixel_index <= 4121)) || ((pixel_index >= 4160) && (pixel_index <= 4162)) || ((pixel_index >= 4209) && (pixel_index <= 4217)) || ((pixel_index >= 4232) && (pixel_index <= 4238)) || ((pixel_index >= 4254) && (pixel_index <= 4259)) || ((pixel_index >= 4306) && (pixel_index <= 4313)) || ((pixel_index >= 4327) && (pixel_index <= 4335)) || ((pixel_index >= 4339) && (pixel_index <= 4341)) || ((pixel_index >= 4348) && (pixel_index <= 4355)) || ((pixel_index >= 4403) && (pixel_index <= 4409)) || ((pixel_index >= 4423) && (pixel_index <= 4439)) || ((pixel_index >= 4443) && (pixel_index <= 4452)) || ((pixel_index >= 4500) && (pixel_index <= 4505)) || ((pixel_index >= 4518) && (pixel_index <= 4548)) || pixel_index == 4570 || ((pixel_index >= 4575) && (pixel_index <= 4577)) || ((pixel_index >= 4583) && (pixel_index <= 4585)) || ((pixel_index >= 4587) && (pixel_index <= 4588)) || ((pixel_index >= 4597) && (pixel_index <= 4601)) || ((pixel_index >= 4613) && (pixel_index <= 4644)) || ((pixel_index >= 4666) && (pixel_index <= 4667)) || ((pixel_index >= 4670) && (pixel_index <= 4675)) || ((pixel_index >= 4677) && (pixel_index <= 4685)) || ((pixel_index >= 4694) && (pixel_index <= 4697)) || ((pixel_index >= 4709) && (pixel_index <= 4740)) || pixel_index == 4757 || ((pixel_index >= 4763) && (pixel_index <= 4781)) || ((pixel_index >= 4791) && (pixel_index <= 4793)) || ((pixel_index >= 4805) && (pixel_index <= 4836)) || pixel_index == 4853 || ((pixel_index >= 4859) && (pixel_index <= 4877)) || ((pixel_index >= 4888) && (pixel_index <= 4889)) || ((pixel_index >= 4901) && (pixel_index <= 4932)) || pixel_index == 4949 || ((pixel_index >= 4955) && (pixel_index <= 4974)) || ((pixel_index >= 4976) && (pixel_index <= 4981)) || pixel_index == 4985 || ((pixel_index >= 4997) && (pixel_index <= 5029)) || pixel_index == 5045 || ((pixel_index >= 5050) && (pixel_index <= 5081)) || ((pixel_index >= 5093) && (pixel_index <= 5125)) || ((pixel_index >= 5141) && (pixel_index <= 5142)) || ((pixel_index >= 5145) && (pixel_index <= 5177)) || ((pixel_index >= 5189) && (pixel_index <= 5221)) || ((pixel_index >= 5237) && (pixel_index <= 5273)) || ((pixel_index >= 5285) && (pixel_index <= 5317)) || ((pixel_index >= 5333) && (pixel_index <= 5369)) || ((pixel_index >= 5381) && (pixel_index <= 5411)) || ((pixel_index >= 5429) && (pixel_index <= 5465)) || ((pixel_index >= 5477) && (pixel_index <= 5507)) || ((pixel_index >= 5525) && (pixel_index <= 5561)) || ((pixel_index >= 5573) && (pixel_index <= 5603)) || ((pixel_index >= 5622) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5700)) || ((pixel_index >= 5718) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5795)) || ((pixel_index >= 5814) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5891)) || ((pixel_index >= 5910) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 5986)) || ((pixel_index >= 6006) && (pixel_index <= 6041)) || ((pixel_index >= 6053) && (pixel_index <= 6082)) || (pixel_index >= 6102) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 3) begin
            if (((pixel_index >= 5) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 377)) || ((pixel_index >= 389) && (pixel_index <= 473)) || ((pixel_index >= 485) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 808)) || ((pixel_index >= 819) && (pixel_index <= 857)) || ((pixel_index >= 869) && (pixel_index <= 903)) || ((pixel_index >= 918) && (pixel_index <= 953)) || ((pixel_index >= 965) && (pixel_index <= 998)) || ((pixel_index >= 1015) && (pixel_index <= 1019)) || ((pixel_index >= 1021) && (pixel_index <= 1049)) || ((pixel_index >= 1061) && (pixel_index <= 1093)) || ((pixel_index >= 1112) && (pixel_index <= 1113)) || ((pixel_index >= 1117) && (pixel_index <= 1145)) || ((pixel_index >= 1157) && (pixel_index <= 1189)) || ((pixel_index >= 1213) && (pixel_index <= 1241)) || ((pixel_index >= 1253) && (pixel_index <= 1285)) || ((pixel_index >= 1309) && (pixel_index <= 1337)) || ((pixel_index >= 1349) && (pixel_index <= 1380)) || ((pixel_index >= 1406) && (pixel_index <= 1433)) || ((pixel_index >= 1445) && (pixel_index <= 1476)) || ((pixel_index >= 1502) && (pixel_index <= 1529)) || ((pixel_index >= 1541) && (pixel_index <= 1572)) || ((pixel_index >= 1599) && (pixel_index <= 1625)) || ((pixel_index >= 1637) && (pixel_index <= 1668)) || ((pixel_index >= 1695) && (pixel_index <= 1721)) || ((pixel_index >= 1733) && (pixel_index <= 1762)) || ((pixel_index >= 1788) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1857)) || ((pixel_index >= 1884) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 1953)) || ((pixel_index >= 1980) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2050)) || ((pixel_index >= 2074) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2147)) || ((pixel_index >= 2170) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2244)) || ((pixel_index >= 2266) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2340)) || ((pixel_index >= 2360) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2436)) || ((pixel_index >= 2455) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2531)) || ((pixel_index >= 2551) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2628)) || ((pixel_index >= 2648) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2725)) || ((pixel_index >= 2743) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2823)) || ((pixel_index >= 2838) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2921)) || ((pixel_index >= 2932) && (pixel_index <= 2969)) || ((pixel_index >= 2981) && (pixel_index <= 2985)) || ((pixel_index >= 2988) && (pixel_index <= 3018)) || ((pixel_index >= 3025) && (pixel_index <= 3065)) || ((pixel_index >= 3077) && (pixel_index <= 3080)) || ((pixel_index >= 3085) && (pixel_index <= 3110)) || ((pixel_index >= 3122) && (pixel_index <= 3161)) || ((pixel_index >= 3173) && (pixel_index <= 3175)) || ((pixel_index >= 3183) && (pixel_index <= 3203)) || ((pixel_index >= 3221) && (pixel_index <= 3257)) || ((pixel_index >= 3269) && (pixel_index <= 3270)) || ((pixel_index >= 3280) && (pixel_index <= 3298)) || ((pixel_index >= 3319) && (pixel_index <= 3338)) || ((pixel_index >= 3340) && (pixel_index <= 3353)) || pixel_index == 3365 || ((pixel_index >= 3378) && (pixel_index <= 3394)) || ((pixel_index >= 3416) && (pixel_index <= 3433)) || ((pixel_index >= 3437) && (pixel_index <= 3449)) || ((pixel_index >= 3475) && (pixel_index <= 3489)) || ((pixel_index >= 3513) && (pixel_index <= 3525)) || ((pixel_index >= 3533) && (pixel_index <= 3545)) || ((pixel_index >= 3572) && (pixel_index <= 3585)) || ((pixel_index >= 3609) && (pixel_index <= 3619)) || ((pixel_index >= 3630) && (pixel_index <= 3641)) || ((pixel_index >= 3670) && (pixel_index <= 3681)) || ((pixel_index >= 3706) && (pixel_index <= 3714)) || ((pixel_index >= 3727) && (pixel_index <= 3737)) || ((pixel_index >= 3774) && (pixel_index <= 3776)) || ((pixel_index >= 3802) && (pixel_index <= 3808)) || ((pixel_index >= 3823) && (pixel_index <= 3833)) || ((pixel_index >= 3920) && (pixel_index <= 3929)) || ((pixel_index >= 4017) && (pixel_index <= 4025)) || ((pixel_index >= 4064) && (pixel_index <= 4066)) || ((pixel_index >= 4114) && (pixel_index <= 4121)) || ((pixel_index >= 4135) && (pixel_index <= 4136)) || ((pixel_index >= 4138) && (pixel_index <= 4140)) || ((pixel_index >= 4158) && (pixel_index <= 4162)) || ((pixel_index >= 4211) && (pixel_index <= 4217)) || ((pixel_index >= 4230) && (pixel_index <= 4237)) || ((pixel_index >= 4252) && (pixel_index <= 4258)) || ((pixel_index >= 4308) && (pixel_index <= 4313)) || ((pixel_index >= 4325) && (pixel_index <= 4334)) || ((pixel_index >= 4337) && (pixel_index <= 4341)) || ((pixel_index >= 4347) && (pixel_index <= 4355)) || pixel_index == 4377 || ((pixel_index >= 4405) && (pixel_index <= 4409)) || ((pixel_index >= 4421) && (pixel_index <= 4438)) || ((pixel_index >= 4441) && (pixel_index <= 4451)) || ((pixel_index >= 4473) && (pixel_index <= 4474)) || ((pixel_index >= 4479) && (pixel_index <= 4481)) || ((pixel_index >= 4487) && (pixel_index <= 4489)) || ((pixel_index >= 4491) && (pixel_index <= 4493)) || ((pixel_index >= 4502) && (pixel_index <= 4505)) || ((pixel_index >= 4517) && (pixel_index <= 4547)) || ((pixel_index >= 4569) && (pixel_index <= 4571)) || ((pixel_index >= 4573) && (pixel_index <= 4579)) || ((pixel_index >= 4581) && (pixel_index <= 4589)) || ((pixel_index >= 4600) && (pixel_index <= 4601)) || ((pixel_index >= 4613) && (pixel_index <= 4643)) || ((pixel_index >= 4665) && (pixel_index <= 4686)) || pixel_index == 4697 || ((pixel_index >= 4709) && (pixel_index <= 4739)) || pixel_index == 4756 || ((pixel_index >= 4762) && (pixel_index <= 4782)) || ((pixel_index >= 4805) && (pixel_index <= 4835)) || pixel_index == 4852 || ((pixel_index >= 4858) && (pixel_index <= 4887)) || ((pixel_index >= 4901) && (pixel_index <= 4931)) || pixel_index == 4948 || ((pixel_index >= 4954) && (pixel_index <= 4985)) || ((pixel_index >= 4997) && (pixel_index <= 5027)) || ((pixel_index >= 5044) && (pixel_index <= 5045)) || ((pixel_index >= 5050) && (pixel_index <= 5081)) || ((pixel_index >= 5093) && (pixel_index <= 5124)) || ((pixel_index >= 5140) && (pixel_index <= 5141)) || ((pixel_index >= 5145) && (pixel_index <= 5177)) || ((pixel_index >= 5189) && (pixel_index <= 5221)) || ((pixel_index >= 5236) && (pixel_index <= 5273)) || ((pixel_index >= 5285) && (pixel_index <= 5316)) || ((pixel_index >= 5332) && (pixel_index <= 5369)) || ((pixel_index >= 5381) && (pixel_index <= 5411)) || ((pixel_index >= 5429) && (pixel_index <= 5465)) || ((pixel_index >= 5477) && (pixel_index <= 5506)) || ((pixel_index >= 5525) && (pixel_index <= 5561)) || ((pixel_index >= 5573) && (pixel_index <= 5603)) || ((pixel_index >= 5622) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5700)) || ((pixel_index >= 5718) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5795)) || ((pixel_index >= 5814) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5890)) || ((pixel_index >= 5910) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 5986)) || ((pixel_index >= 6006) && (pixel_index <= 6041)) || ((pixel_index >= 6053) && (pixel_index <= 6081)) || (pixel_index >= 6102) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 4) begin
            if (((pixel_index >= 5) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 377)) || ((pixel_index >= 389) && (pixel_index <= 473)) || ((pixel_index >= 485) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 857)) || ((pixel_index >= 869) && (pixel_index <= 905)) || ((pixel_index >= 914) && (pixel_index <= 953)) || ((pixel_index >= 965) && (pixel_index <= 999)) || ((pixel_index >= 1014) && (pixel_index <= 1049)) || ((pixel_index >= 1061) && (pixel_index <= 1094)) || ((pixel_index >= 1111) && (pixel_index <= 1145)) || ((pixel_index >= 1157) && (pixel_index <= 1190)) || ((pixel_index >= 1208) && (pixel_index <= 1209)) || ((pixel_index >= 1213) && (pixel_index <= 1241)) || ((pixel_index >= 1253) && (pixel_index <= 1285)) || ((pixel_index >= 1309) && (pixel_index <= 1337)) || ((pixel_index >= 1349) && (pixel_index <= 1381)) || ((pixel_index >= 1405) && (pixel_index <= 1433)) || ((pixel_index >= 1445) && (pixel_index <= 1477)) || ((pixel_index >= 1502) && (pixel_index <= 1529)) || ((pixel_index >= 1541) && (pixel_index <= 1573)) || ((pixel_index >= 1598) && (pixel_index <= 1625)) || ((pixel_index >= 1637) && (pixel_index <= 1669)) || ((pixel_index >= 1694) && (pixel_index <= 1721)) || ((pixel_index >= 1733) && (pixel_index <= 1765)) || ((pixel_index >= 1791) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1859)) || ((pixel_index >= 1884) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 1954)) || ((pixel_index >= 1980) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2049)) || ((pixel_index >= 2076) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2146)) || pixel_index == 2170 || ((pixel_index >= 2172) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2243)) || ((pixel_index >= 2266) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2341)) || ((pixel_index >= 2362) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2437)) || ((pixel_index >= 2456) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2532)) || ((pixel_index >= 2551) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2627)) || ((pixel_index >= 2647) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2724)) || ((pixel_index >= 2744) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2822)) || ((pixel_index >= 2840) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2919)) || ((pixel_index >= 2935) && (pixel_index <= 2969)) || ((pixel_index >= 2981) && (pixel_index <= 2987)) || ((pixel_index >= 2990) && (pixel_index <= 3018)) || ((pixel_index >= 3029) && (pixel_index <= 3065)) || ((pixel_index >= 3077) && (pixel_index <= 3083)) || ((pixel_index >= 3086) && (pixel_index <= 3114)) || ((pixel_index >= 3121) && (pixel_index <= 3161)) || ((pixel_index >= 3173) && (pixel_index <= 3178)) || ((pixel_index >= 3184) && (pixel_index <= 3208)) || ((pixel_index >= 3218) && (pixel_index <= 3257)) || ((pixel_index >= 3269) && (pixel_index <= 3273)) || ((pixel_index >= 3281) && (pixel_index <= 3300)) || ((pixel_index >= 3318) && (pixel_index <= 3339)) || ((pixel_index >= 3341) && (pixel_index <= 3353)) || ((pixel_index >= 3365) && (pixel_index <= 3368)) || ((pixel_index >= 3379) && (pixel_index <= 3395)) || ((pixel_index >= 3416) && (pixel_index <= 3434)) || ((pixel_index >= 3438) && (pixel_index <= 3449)) || ((pixel_index >= 3461) && (pixel_index <= 3463)) || ((pixel_index >= 3476) && (pixel_index <= 3490)) || ((pixel_index >= 3513) && (pixel_index <= 3527)) || ((pixel_index >= 3534) && (pixel_index <= 3545)) || ((pixel_index >= 3557) && (pixel_index <= 3558)) || ((pixel_index >= 3573) && (pixel_index <= 3586)) || ((pixel_index >= 3609) && (pixel_index <= 3621)) || ((pixel_index >= 3631) && (pixel_index <= 3641)) || pixel_index == 3653 || ((pixel_index >= 3670) && (pixel_index <= 3681)) || ((pixel_index >= 3706) && (pixel_index <= 3715)) || ((pixel_index >= 3728) && (pixel_index <= 3737)) || ((pixel_index >= 3768) && (pixel_index <= 3777)) || ((pixel_index >= 3802) && (pixel_index <= 3809)) || ((pixel_index >= 3824) && (pixel_index <= 3833)) || ((pixel_index >= 3871) && (pixel_index <= 3873)) || ((pixel_index >= 3921) && (pixel_index <= 3929)) || ((pixel_index >= 4018) && (pixel_index <= 4025)) || ((pixel_index >= 4115) && (pixel_index <= 4121)) || ((pixel_index >= 4137) && (pixel_index <= 4138)) || pixel_index == 4141 || ((pixel_index >= 4161) && (pixel_index <= 4162)) || ((pixel_index >= 4212) && (pixel_index <= 4217)) || ((pixel_index >= 4232) && (pixel_index <= 4238)) || ((pixel_index >= 4255) && (pixel_index <= 4258)) || ((pixel_index >= 4309) && (pixel_index <= 4313)) || ((pixel_index >= 4328) && (pixel_index <= 4335)) || ((pixel_index >= 4340) && (pixel_index <= 4341)) || ((pixel_index >= 4349) && (pixel_index <= 4354)) || ((pixel_index >= 4406) && (pixel_index <= 4409)) || pixel_index == 4421 || ((pixel_index >= 4423) && (pixel_index <= 4438)) || ((pixel_index >= 4444) && (pixel_index <= 4451)) || ((pixel_index >= 4473) && (pixel_index <= 4475)) || pixel_index == 4481 || ((pixel_index >= 4489) && (pixel_index <= 4490)) || pixel_index == 4493 || ((pixel_index >= 4503) && (pixel_index <= 4505)) || ((pixel_index >= 4517) && (pixel_index <= 4535)) || ((pixel_index >= 4539) && (pixel_index <= 4547)) || ((pixel_index >= 4569) && (pixel_index <= 4572)) || ((pixel_index >= 4575) && (pixel_index <= 4579)) || ((pixel_index >= 4583) && (pixel_index <= 4590)) || ((pixel_index >= 4600) && (pixel_index <= 4601)) || ((pixel_index >= 4613) && (pixel_index <= 4643)) || ((pixel_index >= 4665) && (pixel_index <= 4687)) || pixel_index == 4697 || ((pixel_index >= 4709) && (pixel_index <= 4739)) || ((pixel_index >= 4761) && (pixel_index <= 4783)) || ((pixel_index >= 4805) && (pixel_index <= 4835)) || ((pixel_index >= 4858) && (pixel_index <= 4880)) || ((pixel_index >= 4901) && (pixel_index <= 4931)) || ((pixel_index >= 4954) && (pixel_index <= 4984)) || ((pixel_index >= 4997) && (pixel_index <= 5027)) || ((pixel_index >= 5050) && (pixel_index <= 5081)) || ((pixel_index >= 5093) && (pixel_index <= 5123)) || ((pixel_index >= 5146) && (pixel_index <= 5177)) || ((pixel_index >= 5189) && (pixel_index <= 5221)) || ((pixel_index >= 5237) && (pixel_index <= 5238)) || ((pixel_index >= 5240) && (pixel_index <= 5273)) || ((pixel_index >= 5285) && (pixel_index <= 5317)) || ((pixel_index >= 5333) && (pixel_index <= 5369)) || ((pixel_index >= 5381) && (pixel_index <= 5413)) || ((pixel_index >= 5429) && (pixel_index <= 5465)) || ((pixel_index >= 5477) && (pixel_index <= 5508)) || ((pixel_index >= 5526) && (pixel_index <= 5561)) || ((pixel_index >= 5573) && (pixel_index <= 5604)) || ((pixel_index >= 5623) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5700)) || ((pixel_index >= 5719) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5797)) || ((pixel_index >= 5815) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5892)) || ((pixel_index >= 5911) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 5988)) || ((pixel_index >= 6007) && (pixel_index <= 6041)) || ((pixel_index >= 6053) && (pixel_index <= 6083)) || (pixel_index >= 6103) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 5) begin
            if (((pixel_index >= 5) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 377)) || ((pixel_index >= 389) && (pixel_index <= 473)) || ((pixel_index >= 485) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 809)) || ((pixel_index >= 820) && (pixel_index <= 826)) || ((pixel_index >= 829) && (pixel_index <= 857)) || ((pixel_index >= 869) && (pixel_index <= 903)) || ((pixel_index >= 918) && (pixel_index <= 921)) || ((pixel_index >= 925) && (pixel_index <= 953)) || ((pixel_index >= 965) && (pixel_index <= 998)) || ((pixel_index >= 1015) && (pixel_index <= 1016)) || ((pixel_index >= 1021) && (pixel_index <= 1049)) || ((pixel_index >= 1061) && (pixel_index <= 1094)) || ((pixel_index >= 1118) && (pixel_index <= 1145)) || ((pixel_index >= 1157) && (pixel_index <= 1189)) || ((pixel_index >= 1214) && (pixel_index <= 1241)) || ((pixel_index >= 1253) && (pixel_index <= 1285)) || ((pixel_index >= 1311) && (pixel_index <= 1337)) || ((pixel_index >= 1349) && (pixel_index <= 1381)) || ((pixel_index >= 1408) && (pixel_index <= 1433)) || ((pixel_index >= 1445) && (pixel_index <= 1477)) || ((pixel_index >= 1503) && (pixel_index <= 1529)) || ((pixel_index >= 1541) && (pixel_index <= 1573)) || ((pixel_index >= 1597) && (pixel_index <= 1625)) || ((pixel_index >= 1637) && (pixel_index <= 1669)) || ((pixel_index >= 1693) && (pixel_index <= 1721)) || ((pixel_index >= 1733) && (pixel_index <= 1765)) || ((pixel_index >= 1789) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1859)) || ((pixel_index >= 1882) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 1954)) || ((pixel_index >= 1979) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2050)) || ((pixel_index >= 2075) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2147)) || ((pixel_index >= 2170) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2244)) || ((pixel_index >= 2265) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2342)) || ((pixel_index >= 2360) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2438)) || ((pixel_index >= 2457) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2534)) || ((pixel_index >= 2554) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2629)) || ((pixel_index >= 2649) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2726)) || ((pixel_index >= 2744) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2824)) || ((pixel_index >= 2838) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2896)) || ((pixel_index >= 2898) && (pixel_index <= 2921)) || ((pixel_index >= 2931) && (pixel_index <= 2969)) || ((pixel_index >= 2981) && (pixel_index <= 2991)) || ((pixel_index >= 2995) && (pixel_index <= 3020)) || ((pixel_index >= 3027) && (pixel_index <= 3065)) || ((pixel_index >= 3077) && (pixel_index <= 3086)) || ((pixel_index >= 3092) && (pixel_index <= 3112)) || ((pixel_index >= 3126) && (pixel_index <= 3150)) || ((pixel_index >= 3152) && (pixel_index <= 3161)) || ((pixel_index >= 3173) && (pixel_index <= 3181)) || ((pixel_index >= 3190) && (pixel_index <= 3205)) || ((pixel_index >= 3225) && (pixel_index <= 3246)) || ((pixel_index >= 3249) && (pixel_index <= 3257)) || ((pixel_index >= 3269) && (pixel_index <= 3276)) || ((pixel_index >= 3287) && (pixel_index <= 3300)) || ((pixel_index >= 3322) && (pixel_index <= 3339)) || ((pixel_index >= 3346) && (pixel_index <= 3353)) || ((pixel_index >= 3365) && (pixel_index <= 3371)) || ((pixel_index >= 3384) && (pixel_index <= 3396)) || ((pixel_index >= 3419) && (pixel_index <= 3433)) || ((pixel_index >= 3442) && (pixel_index <= 3449)) || ((pixel_index >= 3461) && (pixel_index <= 3466)) || ((pixel_index >= 3481) && (pixel_index <= 3491)) || ((pixel_index >= 3515) && (pixel_index <= 3527)) || ((pixel_index >= 3539) && (pixel_index <= 3545)) || ((pixel_index >= 3557) && (pixel_index <= 3560)) || ((pixel_index >= 3578) && (pixel_index <= 3587)) || ((pixel_index >= 3612) && (pixel_index <= 3622)) || ((pixel_index >= 3636) && (pixel_index <= 3641)) || ((pixel_index >= 3653) && (pixel_index <= 3655)) || ((pixel_index >= 3676) && (pixel_index <= 3682)) || ((pixel_index >= 3709) && (pixel_index <= 3716)) || ((pixel_index >= 3733) && (pixel_index <= 3737)) || pixel_index == 3749 || ((pixel_index >= 3829) && (pixel_index <= 3833)) || ((pixel_index >= 3926) && (pixel_index <= 3929)) || ((pixel_index >= 4023) && (pixel_index <= 4025)) || ((pixel_index >= 4045) && (pixel_index <= 4046)) || ((pixel_index >= 4048) && (pixel_index <= 4050)) || pixel_index == 4121 || ((pixel_index >= 4140) && (pixel_index <= 4147)) || ((pixel_index >= 4187) && (pixel_index <= 4188)) || ((pixel_index >= 4229) && (pixel_index <= 4230)) || ((pixel_index >= 4235) && (pixel_index <= 4244)) || ((pixel_index >= 4247) && (pixel_index <= 4249)) || ((pixel_index >= 4257) && (pixel_index <= 4259)) || ((pixel_index >= 4283) && (pixel_index <= 4285)) || ((pixel_index >= 4301) && (pixel_index <= 4302)) || ((pixel_index >= 4304) && (pixel_index <= 4305)) || ((pixel_index >= 4325) && (pixel_index <= 4328)) || ((pixel_index >= 4330) && (pixel_index <= 4346)) || ((pixel_index >= 4352) && (pixel_index <= 4356)) || ((pixel_index >= 4379) && (pixel_index <= 4383)) || ((pixel_index >= 4388) && (pixel_index <= 4391)) || ((pixel_index >= 4395) && (pixel_index <= 4402)) || ((pixel_index >= 4421) && (pixel_index <= 4443)) || ((pixel_index >= 4446) && (pixel_index <= 4452)) || ((pixel_index >= 4474) && (pixel_index <= 4480)) || ((pixel_index >= 4482) && (pixel_index <= 4488)) || ((pixel_index >= 4490) && (pixel_index <= 4498)) || ((pixel_index >= 4517) && (pixel_index <= 4548)) || ((pixel_index >= 4570) && (pixel_index <= 4595)) || ((pixel_index >= 4600) && (pixel_index <= 4601)) || ((pixel_index >= 4613) && (pixel_index <= 4644)) || ((pixel_index >= 4666) && (pixel_index <= 4697)) || ((pixel_index >= 4709) && (pixel_index <= 4740)) || ((pixel_index >= 4763) && (pixel_index <= 4793)) || ((pixel_index >= 4805) && (pixel_index <= 4835)) || ((pixel_index >= 4859) && (pixel_index <= 4889)) || ((pixel_index >= 4901) && (pixel_index <= 4932)) || ((pixel_index >= 4955) && (pixel_index <= 4985)) || ((pixel_index >= 4997) && (pixel_index <= 5028)) || ((pixel_index >= 5050) && (pixel_index <= 5081)) || ((pixel_index >= 5093) && (pixel_index <= 5127)) || ((pixel_index >= 5144) && (pixel_index <= 5177)) || ((pixel_index >= 5189) && (pixel_index <= 5223)) || ((pixel_index >= 5240) && (pixel_index <= 5273)) || ((pixel_index >= 5285) && (pixel_index <= 5319)) || ((pixel_index >= 5336) && (pixel_index <= 5369)) || ((pixel_index >= 5381) && (pixel_index <= 5414)) || ((pixel_index >= 5433) && (pixel_index <= 5465)) || ((pixel_index >= 5477) && (pixel_index <= 5510)) || ((pixel_index >= 5530) && (pixel_index <= 5561)) || ((pixel_index >= 5573) && (pixel_index <= 5606)) || ((pixel_index >= 5625) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5702)) || ((pixel_index >= 5721) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5799)) || ((pixel_index >= 5817) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5894)) || ((pixel_index >= 5914) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 5990)) || ((pixel_index >= 6010) && (pixel_index <= 6041)) || ((pixel_index >= 6053) && (pixel_index <= 6086)) || (pixel_index >= 6107) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 6) begin
            if (((pixel_index >= 5) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 377)) || ((pixel_index >= 389) && (pixel_index <= 473)) || ((pixel_index >= 485) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 857)) || ((pixel_index >= 869) && (pixel_index <= 921)) || ((pixel_index >= 923) && (pixel_index <= 953)) || ((pixel_index >= 965) && (pixel_index <= 1006)) || ((pixel_index >= 1011) && (pixel_index <= 1016)) || ((pixel_index >= 1020) && (pixel_index <= 1049)) || ((pixel_index >= 1061) && (pixel_index <= 1096)) || ((pixel_index >= 1109) && (pixel_index <= 1111)) || ((pixel_index >= 1116) && (pixel_index <= 1145)) || ((pixel_index >= 1157) && (pixel_index <= 1191)) || ((pixel_index >= 1213) && (pixel_index <= 1241)) || ((pixel_index >= 1253) && (pixel_index <= 1286)) || ((pixel_index >= 1309) && (pixel_index <= 1337)) || ((pixel_index >= 1349) && (pixel_index <= 1381)) || ((pixel_index >= 1406) && (pixel_index <= 1433)) || ((pixel_index >= 1445) && (pixel_index <= 1477)) || ((pixel_index >= 1503) && (pixel_index <= 1529)) || ((pixel_index >= 1541) && (pixel_index <= 1573)) || ((pixel_index >= 1597) && (pixel_index <= 1625)) || ((pixel_index >= 1637) && (pixel_index <= 1668)) || ((pixel_index >= 1692) && (pixel_index <= 1721)) || ((pixel_index >= 1733) && (pixel_index <= 1764)) || ((pixel_index >= 1788) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1861)) || ((pixel_index >= 1885) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 1957)) || ((pixel_index >= 1977) && (pixel_index <= 1978)) || ((pixel_index >= 1980) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2053)) || ((pixel_index >= 2074) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2148)) || ((pixel_index >= 2171) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2242)) || ((pixel_index >= 2267) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2338)) || ((pixel_index >= 2361) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2434)) || ((pixel_index >= 2457) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2532)) || ((pixel_index >= 2553) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2631)) || ((pixel_index >= 2649) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2726)) || ((pixel_index >= 2746) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2822)) || ((pixel_index >= 2841) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2918)) || ((pixel_index >= 2936) && (pixel_index <= 2969)) || ((pixel_index >= 2981) && (pixel_index <= 3016)) || ((pixel_index >= 3030) && (pixel_index <= 3065)) || ((pixel_index >= 3077) && (pixel_index <= 3113)) || ((pixel_index >= 3123) && (pixel_index <= 3161)) || ((pixel_index >= 3173) && (pixel_index <= 3187)) || ((pixel_index >= 3190) && (pixel_index <= 3212)) || ((pixel_index >= 3219) && (pixel_index <= 3257)) || ((pixel_index >= 3269) && (pixel_index <= 3282)) || ((pixel_index >= 3287) && (pixel_index <= 3307)) || ((pixel_index >= 3319) && (pixel_index <= 3344)) || ((pixel_index >= 3347) && (pixel_index <= 3353)) || ((pixel_index >= 3365) && (pixel_index <= 3377)) || ((pixel_index >= 3385) && (pixel_index <= 3399)) || ((pixel_index >= 3418) && (pixel_index <= 3438)) || ((pixel_index >= 3444) && (pixel_index <= 3449)) || ((pixel_index >= 3461) && (pixel_index <= 3472)) || ((pixel_index >= 3482) && (pixel_index <= 3493)) || ((pixel_index >= 3515) && (pixel_index <= 3532)) || ((pixel_index >= 3540) && (pixel_index <= 3545)) || ((pixel_index >= 3557) && (pixel_index <= 3566)) || ((pixel_index >= 3579) && (pixel_index <= 3589)) || ((pixel_index >= 3611) && (pixel_index <= 3626)) || ((pixel_index >= 3637) && (pixel_index <= 3641)) || ((pixel_index >= 3653) && (pixel_index <= 3661)) || ((pixel_index >= 3676) && (pixel_index <= 3684)) || ((pixel_index >= 3708) && (pixel_index <= 3721)) || ((pixel_index >= 3734) && (pixel_index <= 3737)) || ((pixel_index >= 3749) && (pixel_index <= 3756)) || ((pixel_index >= 3773) && (pixel_index <= 3780)) || ((pixel_index >= 3804) && (pixel_index <= 3815)) || ((pixel_index >= 3830) && (pixel_index <= 3833)) || ((pixel_index >= 3845) && (pixel_index <= 3850)) || ((pixel_index >= 3871) && (pixel_index <= 3875)) || ((pixel_index >= 3901) && (pixel_index <= 3902)) || ((pixel_index >= 3906) && (pixel_index <= 3908)) || ((pixel_index >= 3927) && (pixel_index <= 3929)) || ((pixel_index >= 3941) && (pixel_index <= 3945)) || ((pixel_index >= 3969) && (pixel_index <= 3971)) || ((pixel_index >= 4024) && (pixel_index <= 4025)) || ((pixel_index >= 4037) && (pixel_index <= 4039)) || pixel_index == 4121 || pixel_index == 4133 || ((pixel_index >= 4240) && (pixel_index <= 4241)) || ((pixel_index >= 4244) && (pixel_index <= 4245)) || ((pixel_index >= 4284) && (pixel_index <= 4285)) || ((pixel_index >= 4335) && (pixel_index <= 4342)) || ((pixel_index >= 4380) && (pixel_index <= 4383)) || pixel_index == 4400 || ((pixel_index >= 4402) && (pixel_index <= 4403)) || ((pixel_index >= 4421) && (pixel_index <= 4426)) || ((pixel_index >= 4431) && (pixel_index <= 4439)) || ((pixel_index >= 4442) && (pixel_index <= 4444)) || pixel_index == 4452 || ((pixel_index >= 4475) && (pixel_index <= 4481)) || ((pixel_index >= 4487) && (pixel_index <= 4489)) || ((pixel_index >= 4493) && (pixel_index <= 4496)) || ((pixel_index >= 4498) && (pixel_index <= 4500)) || ((pixel_index >= 4517) && (pixel_index <= 4524)) || ((pixel_index >= 4526) && (pixel_index <= 4541)) || ((pixel_index >= 4546) && (pixel_index <= 4549)) || ((pixel_index >= 4571) && (pixel_index <= 4578)) || ((pixel_index >= 4582) && (pixel_index <= 4586)) || ((pixel_index >= 4589) && (pixel_index <= 4596)) || ((pixel_index >= 4613) && (pixel_index <= 4638)) || ((pixel_index >= 4641) && (pixel_index <= 4645)) || ((pixel_index >= 4667) && (pixel_index <= 4692)) || pixel_index == 4697 || ((pixel_index >= 4709) && (pixel_index <= 4741)) || ((pixel_index >= 4763) && (pixel_index <= 4793)) || ((pixel_index >= 4805) && (pixel_index <= 4836)) || ((pixel_index >= 4859) && (pixel_index <= 4889)) || ((pixel_index >= 4901) && (pixel_index <= 4932)) || ((pixel_index >= 4955) && (pixel_index <= 4985)) || ((pixel_index >= 4997) && (pixel_index <= 5028)) || ((pixel_index >= 5051) && (pixel_index <= 5081)) || ((pixel_index >= 5093) && (pixel_index <= 5125)) || ((pixel_index >= 5147) && (pixel_index <= 5177)) || ((pixel_index >= 5189) && (pixel_index <= 5224)) || ((pixel_index >= 5241) && (pixel_index <= 5273)) || ((pixel_index >= 5285) && (pixel_index <= 5321)) || ((pixel_index >= 5336) && (pixel_index <= 5369)) || ((pixel_index >= 5381) && (pixel_index <= 5417)) || ((pixel_index >= 5432) && (pixel_index <= 5465)) || ((pixel_index >= 5477) && (pixel_index <= 5512)) || ((pixel_index >= 5529) && (pixel_index <= 5561)) || ((pixel_index >= 5573) && (pixel_index <= 5608)) || ((pixel_index >= 5626) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5703)) || ((pixel_index >= 5722) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5799)) || ((pixel_index >= 5818) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5895)) || ((pixel_index >= 5914) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 5991)) || ((pixel_index >= 6010) && (pixel_index <= 6041)) || ((pixel_index >= 6053) && (pixel_index <= 6088)) || (pixel_index >= 6107) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 7) begin
            if (((pixel_index >= 5) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 377)) || ((pixel_index >= 389) && (pixel_index <= 473)) || ((pixel_index >= 485) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 813)) || ((pixel_index >= 820) && (pixel_index <= 826)) || ((pixel_index >= 829) && (pixel_index <= 857)) || ((pixel_index >= 869) && (pixel_index <= 904)) || ((pixel_index >= 919) && (pixel_index <= 920)) || ((pixel_index >= 925) && (pixel_index <= 953)) || ((pixel_index >= 965) && (pixel_index <= 999)) || ((pixel_index >= 1021) && (pixel_index <= 1049)) || ((pixel_index >= 1061) && (pixel_index <= 1094)) || ((pixel_index >= 1118) && (pixel_index <= 1145)) || ((pixel_index >= 1157) && (pixel_index <= 1190)) || ((pixel_index >= 1215) && (pixel_index <= 1241)) || ((pixel_index >= 1253) && (pixel_index <= 1285)) || ((pixel_index >= 1311) && (pixel_index <= 1337)) || ((pixel_index >= 1349) && (pixel_index <= 1381)) || ((pixel_index >= 1408) && (pixel_index <= 1433)) || ((pixel_index >= 1445) && (pixel_index <= 1477)) || ((pixel_index >= 1502) && (pixel_index <= 1529)) || ((pixel_index >= 1541) && (pixel_index <= 1573)) || ((pixel_index >= 1597) && (pixel_index <= 1625)) || ((pixel_index >= 1637) && (pixel_index <= 1669)) || ((pixel_index >= 1694) && (pixel_index <= 1721)) || ((pixel_index >= 1733) && (pixel_index <= 1765)) || pixel_index == 1786 || ((pixel_index >= 1790) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1861)) || ((pixel_index >= 1882) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 1956)) || ((pixel_index >= 1979) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2050)) || ((pixel_index >= 2076) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2146)) || ((pixel_index >= 2171) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2243)) || ((pixel_index >= 2266) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2340)) || ((pixel_index >= 2361) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2439)) || ((pixel_index >= 2458) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2535)) || ((pixel_index >= 2554) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2630)) || ((pixel_index >= 2650) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2726)) || ((pixel_index >= 2746) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2824)) || ((pixel_index >= 2840) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2921)) || ((pixel_index >= 2934) && (pixel_index <= 2969)) || ((pixel_index >= 2981) && (pixel_index <= 2996)) || ((pixel_index >= 2998) && (pixel_index <= 3021)) || ((pixel_index >= 3028) && (pixel_index <= 3058)) || ((pixel_index >= 3060) && (pixel_index <= 3065)) || ((pixel_index >= 3077) && (pixel_index <= 3091)) || ((pixel_index >= 3094) && (pixel_index <= 3116)) || ((pixel_index >= 3125) && (pixel_index <= 3152)) || ((pixel_index >= 3157) && (pixel_index <= 3161)) || ((pixel_index >= 3173) && (pixel_index <= 3186)) || ((pixel_index >= 3192) && (pixel_index <= 3209)) || ((pixel_index >= 3226) && (pixel_index <= 3246)) || ((pixel_index >= 3254) && (pixel_index <= 3257)) || ((pixel_index >= 3269) && (pixel_index <= 3281)) || ((pixel_index >= 3290) && (pixel_index <= 3303)) || ((pixel_index >= 3323) && (pixel_index <= 3340)) || ((pixel_index >= 3350) && (pixel_index <= 3353)) || ((pixel_index >= 3365) && (pixel_index <= 3376)) || ((pixel_index >= 3387) && (pixel_index <= 3398)) || ((pixel_index >= 3420) && (pixel_index <= 3435)) || ((pixel_index >= 3447) && (pixel_index <= 3449)) || ((pixel_index >= 3461) && (pixel_index <= 3471)) || ((pixel_index >= 3484) && (pixel_index <= 3493)) || ((pixel_index >= 3516) && (pixel_index <= 3529)) || ((pixel_index >= 3544) && (pixel_index <= 3545)) || ((pixel_index >= 3557) && (pixel_index <= 3566)) || ((pixel_index >= 3581) && (pixel_index <= 3589)) || ((pixel_index >= 3613) && (pixel_index <= 3623)) || pixel_index == 3641 || ((pixel_index >= 3653) && (pixel_index <= 3660)) || ((pixel_index >= 3679) && (pixel_index <= 3684)) || ((pixel_index >= 3709) && (pixel_index <= 3711)) || pixel_index == 3737 || ((pixel_index >= 3749) && (pixel_index <= 3755)) || ((pixel_index >= 3776) && (pixel_index <= 3780)) || ((pixel_index >= 3845) && (pixel_index <= 3849)) || ((pixel_index >= 3941) && (pixel_index <= 3944)) || ((pixel_index >= 4037) && (pixel_index <= 4038)) || ((pixel_index >= 4092) && (pixel_index <= 4095)) || pixel_index == 4116 || pixel_index == 4133 || ((pixel_index >= 4145) && (pixel_index <= 4146)) || ((pixel_index >= 4148) && (pixel_index <= 4150)) || ((pixel_index >= 4188) && (pixel_index <= 4193)) || ((pixel_index >= 4208) && (pixel_index <= 4209)) || ((pixel_index >= 4211) && (pixel_index <= 4213)) || ((pixel_index >= 4240) && (pixel_index <= 4247)) || ((pixel_index >= 4285) && (pixel_index <= 4291)) || ((pixel_index >= 4296) && (pixel_index <= 4299)) || ((pixel_index >= 4302) && (pixel_index <= 4309)) || ((pixel_index >= 4325) && (pixel_index <= 4331)) || ((pixel_index >= 4335) && (pixel_index <= 4344)) || ((pixel_index >= 4347) && (pixel_index <= 4350)) || ((pixel_index >= 4356) && (pixel_index <= 4357)) || ((pixel_index >= 4380) && (pixel_index <= 4388)) || ((pixel_index >= 4391) && (pixel_index <= 4406)) || ((pixel_index >= 4421) && (pixel_index <= 4428)) || ((pixel_index >= 4430) && (pixel_index <= 4447)) || ((pixel_index >= 4451) && (pixel_index <= 4453)) || ((pixel_index >= 4475) && (pixel_index <= 4505)) || ((pixel_index >= 4517) && (pixel_index <= 4549)) || ((pixel_index >= 4572) && (pixel_index <= 4601)) || ((pixel_index >= 4613) && (pixel_index <= 4645)) || ((pixel_index >= 4668) && (pixel_index <= 4697)) || ((pixel_index >= 4709) && (pixel_index <= 4741)) || ((pixel_index >= 4764) && (pixel_index <= 4793)) || ((pixel_index >= 4805) && (pixel_index <= 4837)) || ((pixel_index >= 4860) && (pixel_index <= 4889)) || ((pixel_index >= 4901) && (pixel_index <= 4933)) || ((pixel_index >= 4956) && (pixel_index <= 4985)) || ((pixel_index >= 4997) && (pixel_index <= 5029)) || ((pixel_index >= 5052) && (pixel_index <= 5081)) || ((pixel_index >= 5093) && (pixel_index <= 5127)) || pixel_index == 5129 || ((pixel_index >= 5147) && (pixel_index <= 5177)) || ((pixel_index >= 5189) && (pixel_index <= 5225)) || ((pixel_index >= 5241) && (pixel_index <= 5273)) || ((pixel_index >= 5285) && (pixel_index <= 5321)) || ((pixel_index >= 5337) && (pixel_index <= 5369)) || ((pixel_index >= 5381) && (pixel_index <= 5417)) || ((pixel_index >= 5433) && (pixel_index <= 5465)) || ((pixel_index >= 5477) && (pixel_index <= 5512)) || ((pixel_index >= 5530) && (pixel_index <= 5561)) || ((pixel_index >= 5573) && (pixel_index <= 5608)) || ((pixel_index >= 5627) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5703)) || ((pixel_index >= 5722) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5799)) || ((pixel_index >= 5818) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5895)) || ((pixel_index >= 5915) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 5992)) || ((pixel_index >= 6011) && (pixel_index <= 6041)) || ((pixel_index >= 6053) && (pixel_index <= 6087)) || (pixel_index >= 6108) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 8) begin
            if (((pixel_index >= 5) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 377)) || ((pixel_index >= 389) && (pixel_index <= 473)) || ((pixel_index >= 485) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 829)) || ((pixel_index >= 831) && (pixel_index <= 857)) || ((pixel_index >= 869) && (pixel_index <= 924)) || ((pixel_index >= 927) && (pixel_index <= 953)) || ((pixel_index >= 965) && (pixel_index <= 1003)) || ((pixel_index >= 1014) && (pixel_index <= 1018)) || ((pixel_index >= 1023) && (pixel_index <= 1049)) || ((pixel_index >= 1061) && (pixel_index <= 1097)) || ((pixel_index >= 1112) && (pixel_index <= 1113)) || ((pixel_index >= 1120) && (pixel_index <= 1145)) || ((pixel_index >= 1157) && (pixel_index <= 1192)) || ((pixel_index >= 1216) && (pixel_index <= 1241)) || ((pixel_index >= 1253) && (pixel_index <= 1287)) || ((pixel_index >= 1313) && (pixel_index <= 1337)) || ((pixel_index >= 1349) && (pixel_index <= 1383)) || ((pixel_index >= 1410) && (pixel_index <= 1433)) || ((pixel_index >= 1445) && (pixel_index <= 1478)) || ((pixel_index >= 1506) && (pixel_index <= 1529)) || ((pixel_index >= 1541) && (pixel_index <= 1574)) || ((pixel_index >= 1600) && (pixel_index <= 1625)) || ((pixel_index >= 1637) && (pixel_index <= 1670)) || ((pixel_index >= 1695) && (pixel_index <= 1721)) || ((pixel_index >= 1733) && (pixel_index <= 1766)) || ((pixel_index >= 1791) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1862)) || ((pixel_index >= 1887) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 1958)) || ((pixel_index >= 1979) && (pixel_index <= 1980)) || ((pixel_index >= 1983) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2053)) || ((pixel_index >= 2076) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2147)) || ((pixel_index >= 2173) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2243)) || ((pixel_index >= 2268) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2340)) || ((pixel_index >= 2364) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2437)) || ((pixel_index >= 2459) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2535)) || ((pixel_index >= 2554) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2632)) || ((pixel_index >= 2651) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2727)) || ((pixel_index >= 2747) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2823)) || ((pixel_index >= 2843) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2919)) || ((pixel_index >= 2938) && (pixel_index <= 2969)) || ((pixel_index >= 2981) && (pixel_index <= 3017)) || ((pixel_index >= 3032) && (pixel_index <= 3065)) || ((pixel_index >= 3077) && (pixel_index <= 3093)) || ((pixel_index >= 3095) && (pixel_index <= 3115)) || ((pixel_index >= 3125) && (pixel_index <= 3155)) || ((pixel_index >= 3157) && (pixel_index <= 3161)) || ((pixel_index >= 3173) && (pixel_index <= 3188)) || ((pixel_index >= 3191) && (pixel_index <= 3214)) || ((pixel_index >= 3221) && (pixel_index <= 3251)) || ((pixel_index >= 3254) && (pixel_index <= 3257)) || ((pixel_index >= 3269) && (pixel_index <= 3283)) || ((pixel_index >= 3289) && (pixel_index <= 3308)) || ((pixel_index >= 3319) && (pixel_index <= 3344)) || ((pixel_index >= 3350) && (pixel_index <= 3353)) || ((pixel_index >= 3365) && (pixel_index <= 3378)) || ((pixel_index >= 3387) && (pixel_index <= 3401)) || ((pixel_index >= 3419) && (pixel_index <= 3438)) || ((pixel_index >= 3447) && (pixel_index <= 3449)) || ((pixel_index >= 3461) && (pixel_index <= 3473)) || ((pixel_index >= 3484) && (pixel_index <= 3495)) || ((pixel_index >= 3516) && (pixel_index <= 3532)) || ((pixel_index >= 3544) && (pixel_index <= 3545)) || ((pixel_index >= 3557) && (pixel_index <= 3567)) || ((pixel_index >= 3581) && (pixel_index <= 3590)) || ((pixel_index >= 3612) && (pixel_index <= 3627)) || pixel_index == 3641 || ((pixel_index >= 3653) && (pixel_index <= 3662)) || ((pixel_index >= 3678) && (pixel_index <= 3686)) || ((pixel_index >= 3709) && (pixel_index <= 3721)) || ((pixel_index >= 3749) && (pixel_index <= 3757)) || ((pixel_index >= 3775) && (pixel_index <= 3781)) || ((pixel_index >= 3805) && (pixel_index <= 3808)) || ((pixel_index >= 3845) && (pixel_index <= 3851)) || ((pixel_index >= 3873) && (pixel_index <= 3877)) || ((pixel_index >= 3941) && (pixel_index <= 3945)) || ((pixel_index >= 4037) && (pixel_index <= 4039)) || ((pixel_index >= 4133) && (pixel_index <= 4134)) || pixel_index == 4146 || ((pixel_index >= 4190) && (pixel_index <= 4191)) || ((pixel_index >= 4241) && (pixel_index <= 4243)) || ((pixel_index >= 4245) && (pixel_index <= 4247)) || ((pixel_index >= 4285) && (pixel_index <= 4289)) || ((pixel_index >= 4305) && (pixel_index <= 4306)) || ((pixel_index >= 4308) && (pixel_index <= 4310)) || ((pixel_index >= 4326) && (pixel_index <= 4330)) || ((pixel_index >= 4336) && (pixel_index <= 4344)) || ((pixel_index >= 4381) && (pixel_index <= 4387)) || ((pixel_index >= 4393) && (pixel_index <= 4395)) || ((pixel_index >= 4399) && (pixel_index <= 4406)) || ((pixel_index >= 4421) && (pixel_index <= 4428)) || ((pixel_index >= 4431) && (pixel_index <= 4441)) || ((pixel_index >= 4443) && (pixel_index <= 4447)) || pixel_index == 4453 || ((pixel_index >= 4477) && (pixel_index <= 4485)) || ((pixel_index >= 4488) && (pixel_index <= 4493)) || ((pixel_index >= 4495) && (pixel_index <= 4503)) || ((pixel_index >= 4517) && (pixel_index <= 4544)) || ((pixel_index >= 4547) && (pixel_index <= 4550)) || ((pixel_index >= 4572) && (pixel_index <= 4601)) || ((pixel_index >= 4613) && (pixel_index <= 4646)) || ((pixel_index >= 4668) && (pixel_index <= 4697)) || ((pixel_index >= 4709) && (pixel_index <= 4742)) || ((pixel_index >= 4764) && (pixel_index <= 4793)) || ((pixel_index >= 4805) && (pixel_index <= 4838)) || ((pixel_index >= 4860) && (pixel_index <= 4889)) || ((pixel_index >= 4901) && (pixel_index <= 4934)) || ((pixel_index >= 4957) && (pixel_index <= 4985)) || ((pixel_index >= 4997) && (pixel_index <= 5029)) || ((pixel_index >= 5053) && (pixel_index <= 5081)) || ((pixel_index >= 5093) && (pixel_index <= 5126)) || ((pixel_index >= 5148) && (pixel_index <= 5177)) || ((pixel_index >= 5189) && (pixel_index <= 5223)) || ((pixel_index >= 5244) && (pixel_index <= 5273)) || ((pixel_index >= 5285) && (pixel_index <= 5322)) || ((pixel_index >= 5339) && (pixel_index <= 5369)) || ((pixel_index >= 5381) && (pixel_index <= 5417)) || ((pixel_index >= 5433) && (pixel_index <= 5465)) || ((pixel_index >= 5477) && (pixel_index <= 5513)) || ((pixel_index >= 5529) && (pixel_index <= 5561)) || ((pixel_index >= 5573) && (pixel_index <= 5608)) || ((pixel_index >= 5626) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5704)) || ((pixel_index >= 5722) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5799)) || ((pixel_index >= 5818) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5895)) || ((pixel_index >= 5914) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 5991)) || ((pixel_index >= 6010) && (pixel_index <= 6041)) || ((pixel_index >= 6053) && (pixel_index <= 6088)) || (pixel_index >= 6107) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 9) begin
            if (((pixel_index >= 5) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 377)) || ((pixel_index >= 389) && (pixel_index <= 473)) || ((pixel_index >= 485) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 811)) || ((pixel_index >= 822) && (pixel_index <= 831)) || ((pixel_index >= 834) && (pixel_index <= 857)) || ((pixel_index >= 869) && (pixel_index <= 905)) || ((pixel_index >= 921) && (pixel_index <= 925)) || ((pixel_index >= 930) && (pixel_index <= 953)) || ((pixel_index >= 965) && (pixel_index <= 1000)) || ((pixel_index >= 1018) && (pixel_index <= 1020)) || ((pixel_index >= 1026) && (pixel_index <= 1049)) || ((pixel_index >= 1061) && (pixel_index <= 1095)) || ((pixel_index >= 1122) && (pixel_index <= 1145)) || ((pixel_index >= 1157) && (pixel_index <= 1191)) || ((pixel_index >= 1219) && (pixel_index <= 1241)) || ((pixel_index >= 1253) && (pixel_index <= 1287)) || ((pixel_index >= 1315) && (pixel_index <= 1337)) || ((pixel_index >= 1349) && (pixel_index <= 1382)) || ((pixel_index >= 1412) && (pixel_index <= 1433)) || ((pixel_index >= 1445) && (pixel_index <= 1478)) || ((pixel_index >= 1509) && (pixel_index <= 1529)) || ((pixel_index >= 1541) && (pixel_index <= 1574)) || ((pixel_index >= 1605) && (pixel_index <= 1625)) || ((pixel_index >= 1637) && (pixel_index <= 1670)) || ((pixel_index >= 1698) && (pixel_index <= 1721)) || ((pixel_index >= 1733) && (pixel_index <= 1766)) || ((pixel_index >= 1794) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1861)) || ((pixel_index >= 1890) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 1955)) || ((pixel_index >= 1980) && (pixel_index <= 1981)) || ((pixel_index >= 1985) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2050)) || ((pixel_index >= 2077) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2146)) || ((pixel_index >= 2173) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2243)) || ((pixel_index >= 2269) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2341)) || ((pixel_index >= 2364) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2439)) || ((pixel_index >= 2460) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2535)) || ((pixel_index >= 2555) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2631)) || ((pixel_index >= 2651) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2726)) || ((pixel_index >= 2748) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2823)) || ((pixel_index >= 2844) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2900)) || ((pixel_index >= 2903) && (pixel_index <= 2919)) || ((pixel_index >= 2940) && (pixel_index <= 2969)) || ((pixel_index >= 2981) && (pixel_index <= 2995)) || ((pixel_index >= 2999) && (pixel_index <= 3018)) || ((pixel_index >= 3033) && (pixel_index <= 3065)) || ((pixel_index >= 3077) && (pixel_index <= 3091)) || ((pixel_index >= 3096) && (pixel_index <= 3117)) || ((pixel_index >= 3125) && (pixel_index <= 3126)) || ((pixel_index >= 3128) && (pixel_index <= 3161)) || ((pixel_index >= 3173) && (pixel_index <= 3186)) || ((pixel_index >= 3193) && (pixel_index <= 3213)) || ((pixel_index >= 3221) && (pixel_index <= 3257)) || ((pixel_index >= 3269) && (pixel_index <= 3281)) || ((pixel_index >= 3291) && (pixel_index <= 3305)) || ((pixel_index >= 3318) && (pixel_index <= 3353)) || ((pixel_index >= 3365) && (pixel_index <= 3376)) || ((pixel_index >= 3387) && (pixel_index <= 3398)) || ((pixel_index >= 3417) && (pixel_index <= 3446)) || pixel_index == 3449 || ((pixel_index >= 3461) && (pixel_index <= 3471)) || ((pixel_index >= 3484) && (pixel_index <= 3493)) || ((pixel_index >= 3516) && (pixel_index <= 3540)) || ((pixel_index >= 3557) && (pixel_index <= 3565)) || ((pixel_index >= 3581) && (pixel_index <= 3588)) || ((pixel_index >= 3613) && (pixel_index <= 3633)) || ((pixel_index >= 3653) && (pixel_index <= 3660)) || ((pixel_index >= 3678) && (pixel_index <= 3684)) || ((pixel_index >= 3709) && (pixel_index <= 3727)) || ((pixel_index >= 3749) && (pixel_index <= 3754)) || ((pixel_index >= 3775) && (pixel_index <= 3779)) || ((pixel_index >= 3806) && (pixel_index <= 3822)) || ((pixel_index >= 3845) && (pixel_index <= 3849)) || pixel_index == 3874 || ((pixel_index >= 3902) && (pixel_index <= 3916)) || ((pixel_index >= 3941) && (pixel_index <= 3944)) || ((pixel_index >= 3998) && (pixel_index <= 4000)) || ((pixel_index >= 4005) && (pixel_index <= 4009)) || ((pixel_index >= 4037) && (pixel_index <= 4040)) || pixel_index == 4042 || ((pixel_index >= 4049) && (pixel_index <= 4050)) || ((pixel_index >= 4052) && (pixel_index <= 4053)) || ((pixel_index >= 4133) && (pixel_index <= 4140)) || ((pixel_index >= 4145) && (pixel_index <= 4150)) || ((pixel_index >= 4229) && (pixel_index <= 4238)) || ((pixel_index >= 4240) && (pixel_index <= 4247)) || ((pixel_index >= 4325) && (pixel_index <= 4349)) || pixel_index == 4382 || ((pixel_index >= 4421) && (pixel_index <= 4446)) || ((pixel_index >= 4477) && (pixel_index <= 4480)) || ((pixel_index >= 4517) && (pixel_index <= 4542)) || ((pixel_index >= 4545) && (pixel_index <= 4547)) || ((pixel_index >= 4573) && (pixel_index <= 4578)) || ((pixel_index >= 4613) && (pixel_index <= 4643)) || ((pixel_index >= 4669) && (pixel_index <= 4676)) || ((pixel_index >= 4683) && (pixel_index <= 4684)) || ((pixel_index >= 4692) && (pixel_index <= 4694)) || pixel_index == 4697 || ((pixel_index >= 4709) && (pixel_index <= 4738)) || ((pixel_index >= 4764) && (pixel_index <= 4773)) || ((pixel_index >= 4777) && (pixel_index <= 4782)) || ((pixel_index >= 4786) && (pixel_index <= 4790)) || ((pixel_index >= 4792) && (pixel_index <= 4793)) || ((pixel_index >= 4805) && (pixel_index <= 4834)) || ((pixel_index >= 4859) && (pixel_index <= 4889)) || ((pixel_index >= 4901) && (pixel_index <= 4930)) || ((pixel_index >= 4955) && (pixel_index <= 4985)) || ((pixel_index >= 4997) && (pixel_index <= 5026)) || ((pixel_index >= 5051) && (pixel_index <= 5081)) || ((pixel_index >= 5093) && (pixel_index <= 5122)) || ((pixel_index >= 5147) && (pixel_index <= 5177)) || ((pixel_index >= 5189) && (pixel_index <= 5218)) || ((pixel_index >= 5243) && (pixel_index <= 5273)) || ((pixel_index >= 5285) && (pixel_index <= 5315)) || ((pixel_index >= 5339) && (pixel_index <= 5369)) || ((pixel_index >= 5381) && (pixel_index <= 5415)) || ((pixel_index >= 5435) && (pixel_index <= 5465)) || ((pixel_index >= 5477) && (pixel_index <= 5510)) || ((pixel_index >= 5529) && (pixel_index <= 5561)) || ((pixel_index >= 5573) && (pixel_index <= 5606)) || ((pixel_index >= 5623) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5702)) || ((pixel_index >= 5719) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5797)) || ((pixel_index >= 5816) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5893)) || ((pixel_index >= 5913) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 5988)) || ((pixel_index >= 6009) && (pixel_index <= 6041)) || ((pixel_index >= 6053) && (pixel_index <= 6084)) || (pixel_index >= 6105) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 10) begin
            if (((pixel_index >= 5) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 377)) || ((pixel_index >= 389) && (pixel_index <= 473)) || ((pixel_index >= 485) && (pixel_index <= 527)) || ((pixel_index >= 533) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 618)) || ((pixel_index >= 633) && (pixel_index <= 641)) || ((pixel_index >= 647) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 713)) || ((pixel_index >= 731) && (pixel_index <= 735)) || ((pixel_index >= 743) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 808)) || ((pixel_index >= 828) && (pixel_index <= 829)) || ((pixel_index >= 839) && (pixel_index <= 857)) || ((pixel_index >= 869) && (pixel_index <= 904)) || ((pixel_index >= 935) && (pixel_index <= 953)) || ((pixel_index >= 965) && (pixel_index <= 999)) || ((pixel_index >= 1031) && (pixel_index <= 1049)) || ((pixel_index >= 1061) && (pixel_index <= 1095)) || ((pixel_index >= 1128) && (pixel_index <= 1145)) || ((pixel_index >= 1157) && (pixel_index <= 1191)) || ((pixel_index >= 1224) && (pixel_index <= 1241)) || ((pixel_index >= 1253) && (pixel_index <= 1286)) || ((pixel_index >= 1321) && (pixel_index <= 1337)) || ((pixel_index >= 1349) && (pixel_index <= 1382)) || ((pixel_index >= 1417) && (pixel_index <= 1433)) || ((pixel_index >= 1445) && (pixel_index <= 1478)) || ((pixel_index >= 1514) && (pixel_index <= 1529)) || ((pixel_index >= 1541) && (pixel_index <= 1571)) || ((pixel_index >= 1606) && (pixel_index <= 1625)) || ((pixel_index >= 1637) && (pixel_index <= 1666)) || ((pixel_index >= 1703) && (pixel_index <= 1721)) || ((pixel_index >= 1733) && (pixel_index <= 1761)) || ((pixel_index >= 1798) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1857)) || ((pixel_index >= 1885) && (pixel_index <= 1886)) || ((pixel_index >= 1894) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 1954)) || ((pixel_index >= 1981) && (pixel_index <= 1985)) || ((pixel_index >= 1989) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2052)) || ((pixel_index >= 2077) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2149)) || ((pixel_index >= 2174) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2246)) || ((pixel_index >= 2269) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2343)) || ((pixel_index >= 2365) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2439)) || ((pixel_index >= 2461) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2535)) || ((pixel_index >= 2557) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2617)) || ((pixel_index >= 2619) && (pixel_index <= 2631)) || ((pixel_index >= 2653) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2713)) || ((pixel_index >= 2716) && (pixel_index <= 2727)) || ((pixel_index >= 2749) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2808)) || ((pixel_index >= 2812) && (pixel_index <= 2824)) || ((pixel_index >= 2845) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2903)) || ((pixel_index >= 2908) && (pixel_index <= 2921)) || ((pixel_index >= 2941) && (pixel_index <= 2969)) || ((pixel_index >= 2981) && (pixel_index <= 2998)) || ((pixel_index >= 3005) && (pixel_index <= 3019)) || pixel_index == 3021 || ((pixel_index >= 3034) && (pixel_index <= 3065)) || ((pixel_index >= 3077) && (pixel_index <= 3093)) || ((pixel_index >= 3102) && (pixel_index <= 3117)) || pixel_index == 3127 || ((pixel_index >= 3130) && (pixel_index <= 3161)) || ((pixel_index >= 3173) && (pixel_index <= 3188)) || ((pixel_index >= 3198) && (pixel_index <= 3213)) || ((pixel_index >= 3221) && (pixel_index <= 3257)) || ((pixel_index >= 3269) && (pixel_index <= 3283)) || ((pixel_index >= 3295) && (pixel_index <= 3302)) || ((pixel_index >= 3318) && (pixel_index <= 3353)) || ((pixel_index >= 3365) && (pixel_index <= 3378)) || ((pixel_index >= 3392) && (pixel_index <= 3398)) || ((pixel_index >= 3416) && (pixel_index <= 3449)) || ((pixel_index >= 3461) && (pixel_index <= 3473)) || ((pixel_index >= 3488) && (pixel_index <= 3493)) || ((pixel_index >= 3514) && (pixel_index <= 3545)) || ((pixel_index >= 3557) && (pixel_index <= 3567)) || ((pixel_index >= 3585) && (pixel_index <= 3588)) || ((pixel_index >= 3612) && (pixel_index <= 3641)) || ((pixel_index >= 3653) && (pixel_index <= 3663)) || ((pixel_index >= 3682) && (pixel_index <= 3683)) || ((pixel_index >= 3709) && (pixel_index <= 3735)) || ((pixel_index >= 3749) && (pixel_index <= 3761)) || ((pixel_index >= 3805) && (pixel_index <= 3828)) || ((pixel_index >= 3845) && (pixel_index <= 3858)) || pixel_index == 3862 || pixel_index == 3864 || ((pixel_index >= 3901) && (pixel_index <= 3922)) || ((pixel_index >= 3941) && (pixel_index <= 3955)) || ((pixel_index >= 3957) && (pixel_index <= 3960)) || ((pixel_index >= 3997) && (pixel_index <= 4016)) || ((pixel_index >= 4037) && (pixel_index <= 4057)) || ((pixel_index >= 4093) && (pixel_index <= 4110)) || ((pixel_index >= 4133) && (pixel_index <= 4153)) || ((pixel_index >= 4190) && (pixel_index <= 4193)) || ((pixel_index >= 4196) && (pixel_index <= 4204)) || ((pixel_index >= 4229) && (pixel_index <= 4248)) || ((pixel_index >= 4325) && (pixel_index <= 4344)) || ((pixel_index >= 4421) && (pixel_index <= 4441)) || ((pixel_index >= 4517) && (pixel_index <= 4539)) || pixel_index == 4573 || ((pixel_index >= 4613) && (pixel_index <= 4636)) || ((pixel_index >= 4668) && (pixel_index <= 4671)) || ((pixel_index >= 4709) && (pixel_index <= 4734)) || ((pixel_index >= 4763) && (pixel_index <= 4769)) || ((pixel_index >= 4805) && (pixel_index <= 4830)) || ((pixel_index >= 4859) && (pixel_index <= 4867)) || ((pixel_index >= 4901) && (pixel_index <= 4926)) || ((pixel_index >= 4955) && (pixel_index <= 4964)) || ((pixel_index >= 4997) && (pixel_index <= 5022)) || ((pixel_index >= 5048) && (pixel_index <= 5061)) || ((pixel_index >= 5067) && (pixel_index <= 5069)) || ((pixel_index >= 5093) && (pixel_index <= 5118)) || ((pixel_index >= 5144) && (pixel_index <= 5159)) || ((pixel_index >= 5162) && (pixel_index <= 5167)) || ((pixel_index >= 5173) && (pixel_index <= 5177)) || ((pixel_index >= 5189) && (pixel_index <= 5214)) || ((pixel_index >= 5240) && (pixel_index <= 5264)) || ((pixel_index >= 5267) && (pixel_index <= 5273)) || ((pixel_index >= 5285) && (pixel_index <= 5311)) || ((pixel_index >= 5336) && (pixel_index <= 5369)) || ((pixel_index >= 5381) && (pixel_index <= 5411)) || ((pixel_index >= 5431) && (pixel_index <= 5465)) || ((pixel_index >= 5477) && (pixel_index <= 5507)) || ((pixel_index >= 5527) && (pixel_index <= 5561)) || ((pixel_index >= 5573) && (pixel_index <= 5603)) || ((pixel_index >= 5623) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5699)) || ((pixel_index >= 5718) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5795)) || ((pixel_index >= 5813) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5890)) || ((pixel_index >= 5909) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 5985)) || ((pixel_index >= 6005) && (pixel_index <= 6041)) || ((pixel_index >= 6053) && (pixel_index <= 6081)) || (pixel_index >= 6102) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 11) begin
            if (((pixel_index >= 5) && (pixel_index <= 47)) || ((pixel_index >= 60) && (pixel_index <= 63)) || ((pixel_index >= 76) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 140)) || pixel_index == 158 || ((pixel_index >= 172) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 235)) || ((pixel_index >= 268) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 330)) || ((pixel_index >= 364) && (pixel_index <= 377)) || ((pixel_index >= 389) && (pixel_index <= 425)) || ((pixel_index >= 460) && (pixel_index <= 473)) || ((pixel_index >= 485) && (pixel_index <= 521)) || ((pixel_index >= 557) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 617)) || ((pixel_index >= 653) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 712)) || ((pixel_index >= 750) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 808)) || ((pixel_index >= 846) && (pixel_index <= 857)) || ((pixel_index >= 869) && (pixel_index <= 904)) || ((pixel_index >= 942) && (pixel_index <= 953)) || ((pixel_index >= 965) && (pixel_index <= 1000)) || ((pixel_index >= 1035) && (pixel_index <= 1049)) || ((pixel_index >= 1061) && (pixel_index <= 1094)) || ((pixel_index >= 1132) && (pixel_index <= 1145)) || ((pixel_index >= 1157) && (pixel_index <= 1189)) || ((pixel_index >= 1228) && (pixel_index <= 1241)) || ((pixel_index >= 1253) && (pixel_index <= 1283)) || ((pixel_index >= 1323) && (pixel_index <= 1337)) || ((pixel_index >= 1349) && (pixel_index <= 1376)) || ((pixel_index >= 1418) && (pixel_index <= 1433)) || ((pixel_index >= 1445) && (pixel_index <= 1472)) || ((pixel_index >= 1505) && (pixel_index <= 1506)) || ((pixel_index >= 1513) && (pixel_index <= 1529)) || ((pixel_index >= 1541) && (pixel_index <= 1569)) || pixel_index == 1571 || ((pixel_index >= 1601) && (pixel_index <= 1605)) || ((pixel_index >= 1607) && (pixel_index <= 1625)) || ((pixel_index >= 1637) && (pixel_index <= 1670)) || ((pixel_index >= 1697) && (pixel_index <= 1721)) || ((pixel_index >= 1733) && (pixel_index <= 1766)) || ((pixel_index >= 1794) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1863)) || ((pixel_index >= 1890) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 1960)) || ((pixel_index >= 1987) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2056)) || ((pixel_index >= 2083) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2154)) || ((pixel_index >= 2179) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2250)) || ((pixel_index >= 2275) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2346)) || ((pixel_index >= 2368) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2442)) || ((pixel_index >= 2464) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2537)) || ((pixel_index >= 2560) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2633)) || ((pixel_index >= 2657) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2728)) || pixel_index == 2734 || ((pixel_index >= 2752) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2824)) || ((pixel_index >= 2830) && (pixel_index <= 2833)) || ((pixel_index >= 2846) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2919)) || ((pixel_index >= 2926) && (pixel_index <= 2929)) || ((pixel_index >= 2937) && (pixel_index <= 2969)) || ((pixel_index >= 2981) && (pixel_index <= 3015)) || ((pixel_index >= 3033) && (pixel_index <= 3065)) || ((pixel_index >= 3077) && (pixel_index <= 3110)) || ((pixel_index >= 3130) && (pixel_index <= 3161)) || ((pixel_index >= 3173) && (pixel_index <= 3206)) || ((pixel_index >= 3228) && (pixel_index <= 3257)) || ((pixel_index >= 3269) && (pixel_index <= 3301)) || ((pixel_index >= 3325) && (pixel_index <= 3353)) || ((pixel_index >= 3365) && (pixel_index <= 3398)) || ((pixel_index >= 3422) && (pixel_index <= 3449)) || ((pixel_index >= 3461) && (pixel_index <= 3494)) || ((pixel_index >= 3519) && (pixel_index <= 3545)) || ((pixel_index >= 3557) && (pixel_index <= 3590)) || ((pixel_index >= 3616) && (pixel_index <= 3641)) || ((pixel_index >= 3653) && (pixel_index <= 3668)) || pixel_index == 3682 || ((pixel_index >= 3684) && (pixel_index <= 3686)) || ((pixel_index >= 3712) && (pixel_index <= 3737)) || ((pixel_index >= 3749) && (pixel_index <= 3764)) || ((pixel_index >= 3808) && (pixel_index <= 3833)) || ((pixel_index >= 3845) && (pixel_index <= 3860)) || ((pixel_index >= 3904) && (pixel_index <= 3929)) || ((pixel_index >= 3941) && (pixel_index <= 3956)) || ((pixel_index >= 4000) && (pixel_index <= 4023)) || ((pixel_index >= 4037) && (pixel_index <= 4053)) || ((pixel_index >= 4097) && (pixel_index <= 4118)) || ((pixel_index >= 4133) && (pixel_index <= 4146)) || ((pixel_index >= 4196) && (pixel_index <= 4212)) || ((pixel_index >= 4229) && (pixel_index <= 4243)) || pixel_index == 4294 || ((pixel_index >= 4301) && (pixel_index <= 4305)) || ((pixel_index >= 4325) && (pixel_index <= 4340)) || ((pixel_index >= 4421) && (pixel_index <= 4438)) || ((pixel_index >= 4517) && (pixel_index <= 4535)) || ((pixel_index >= 4541) && (pixel_index <= 4542)) || ((pixel_index >= 4575) && (pixel_index <= 4578)) || ((pixel_index >= 4613) && (pixel_index <= 4639)) || ((pixel_index >= 4670) && (pixel_index <= 4676)) || ((pixel_index >= 4709) && (pixel_index <= 4735)) || ((pixel_index >= 4763) && (pixel_index <= 4773)) || ((pixel_index >= 4805) && (pixel_index <= 4832)) || ((pixel_index >= 4859) && (pixel_index <= 4871)) || ((pixel_index >= 4901) && (pixel_index <= 4928)) || ((pixel_index >= 4955) && (pixel_index <= 4968)) || ((pixel_index >= 4997) && (pixel_index <= 5025)) || ((pixel_index >= 5049) && (pixel_index <= 5065)) || ((pixel_index >= 5093) && (pixel_index <= 5121)) || ((pixel_index >= 5145) && (pixel_index <= 5162)) || ((pixel_index >= 5189) && (pixel_index <= 5218)) || ((pixel_index >= 5241) && (pixel_index <= 5260)) || ((pixel_index >= 5268) && (pixel_index <= 5269)) || ((pixel_index >= 5285) && (pixel_index <= 5316)) || ((pixel_index >= 5337) && (pixel_index <= 5357)) || ((pixel_index >= 5362) && (pixel_index <= 5367)) || ((pixel_index >= 5381) && (pixel_index <= 5414)) || ((pixel_index >= 5432) && (pixel_index <= 5454)) || ((pixel_index >= 5457) && (pixel_index <= 5464)) || ((pixel_index >= 5477) && (pixel_index <= 5510)) || ((pixel_index >= 5528) && (pixel_index <= 5561)) || ((pixel_index >= 5573) && (pixel_index <= 5606)) || ((pixel_index >= 5624) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5702)) || ((pixel_index >= 5720) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5797)) || ((pixel_index >= 5816) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5893)) || ((pixel_index >= 5912) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 5988)) || ((pixel_index >= 6009) && (pixel_index <= 6041)) || ((pixel_index >= 6053) && (pixel_index <= 6083)) || (pixel_index >= 6106) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 12) begin
            if (((pixel_index >= 5) && (pixel_index <= 62)) || ((pixel_index >= 75) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 157)) || ((pixel_index >= 172) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 248)) || ((pixel_index >= 268) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 341)) || ((pixel_index >= 364) && (pixel_index <= 377)) || ((pixel_index >= 389) && (pixel_index <= 435)) || ((pixel_index >= 460) && (pixel_index <= 473)) || ((pixel_index >= 485) && (pixel_index <= 530)) || ((pixel_index >= 554) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 625)) || ((pixel_index >= 650) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 720)) || ((pixel_index >= 750) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 816)) || ((pixel_index >= 846) && (pixel_index <= 857)) || ((pixel_index >= 869) && (pixel_index <= 911)) || ((pixel_index >= 941) && (pixel_index <= 953)) || ((pixel_index >= 965) && (pixel_index <= 1007)) || ((pixel_index >= 1036) && (pixel_index <= 1049)) || ((pixel_index >= 1061) && (pixel_index <= 1103)) || ((pixel_index >= 1131) && (pixel_index <= 1145)) || ((pixel_index >= 1157) && (pixel_index <= 1199)) || ((pixel_index >= 1226) && (pixel_index <= 1241)) || ((pixel_index >= 1253) && (pixel_index <= 1294)) || ((pixel_index >= 1322) && (pixel_index <= 1337)) || ((pixel_index >= 1349) && (pixel_index <= 1390)) || ((pixel_index >= 1418) && (pixel_index <= 1433)) || ((pixel_index >= 1445) && (pixel_index <= 1484)) || ((pixel_index >= 1513) && (pixel_index <= 1529)) || ((pixel_index >= 1541) && (pixel_index <= 1578)) || ((pixel_index >= 1609) && (pixel_index <= 1625)) || ((pixel_index >= 1637) && (pixel_index <= 1672)) || ((pixel_index >= 1705) && (pixel_index <= 1721)) || ((pixel_index >= 1733) && (pixel_index <= 1768)) || ((pixel_index >= 1801) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1865)) || ((pixel_index >= 1898) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 1965)) || ((pixel_index >= 1994) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2062)) || ((pixel_index >= 2091) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2159)) || ((pixel_index >= 2189) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2257)) || pixel_index == 2281 || ((pixel_index >= 2285) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2354)) || ((pixel_index >= 2377) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2450)) || ((pixel_index >= 2473) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2547)) || ((pixel_index >= 2570) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2643)) || ((pixel_index >= 2666) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2739)) || ((pixel_index >= 2761) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2836)) || pixel_index == 2854 || ((pixel_index >= 2857) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2934)) || ((pixel_index >= 2937) && (pixel_index <= 2938)) || ((pixel_index >= 2947) && (pixel_index <= 2950)) || ((pixel_index >= 2954) && (pixel_index <= 2969)) || ((pixel_index >= 2981) && (pixel_index <= 3033)) || ((pixel_index >= 3042) && (pixel_index <= 3045)) || ((pixel_index >= 3050) && (pixel_index <= 3065)) || ((pixel_index >= 3077) && (pixel_index <= 3129)) || ((pixel_index >= 3138) && (pixel_index <= 3141)) || ((pixel_index >= 3146) && (pixel_index <= 3161)) || ((pixel_index >= 3173) && (pixel_index <= 3223)) || ((pixel_index >= 3234) && (pixel_index <= 3237)) || ((pixel_index >= 3243) && (pixel_index <= 3257)) || ((pixel_index >= 3269) && (pixel_index <= 3318)) || ((pixel_index >= 3331) && (pixel_index <= 3333)) || ((pixel_index >= 3339) && (pixel_index <= 3353)) || ((pixel_index >= 3365) && (pixel_index <= 3413)) || ((pixel_index >= 3427) && (pixel_index <= 3429)) || ((pixel_index >= 3436) && (pixel_index <= 3449)) || ((pixel_index >= 3461) && (pixel_index <= 3509)) || ((pixel_index >= 3524) && (pixel_index <= 3525)) || ((pixel_index >= 3532) && (pixel_index <= 3545)) || ((pixel_index >= 3557) && (pixel_index <= 3576)) || ((pixel_index >= 3588) && (pixel_index <= 3604)) || ((pixel_index >= 3629) && (pixel_index <= 3641)) || ((pixel_index >= 3653) && (pixel_index <= 3672)) || ((pixel_index >= 3687) && (pixel_index <= 3698)) || ((pixel_index >= 3724) && (pixel_index <= 3737)) || ((pixel_index >= 3749) && (pixel_index <= 3768)) || ((pixel_index >= 3785) && (pixel_index <= 3793)) || ((pixel_index >= 3820) && (pixel_index <= 3833)) || ((pixel_index >= 3845) && (pixel_index <= 3865)) || ((pixel_index >= 3883) && (pixel_index <= 3889)) || ((pixel_index >= 3915) && (pixel_index <= 3929)) || ((pixel_index >= 3941) && (pixel_index <= 3961)) || ((pixel_index >= 3979) && (pixel_index <= 3985)) || ((pixel_index >= 4008) && (pixel_index <= 4025)) || ((pixel_index >= 4037) && (pixel_index <= 4056)) || ((pixel_index >= 4076) && (pixel_index <= 4080)) || ((pixel_index >= 4104) && (pixel_index <= 4121)) || ((pixel_index >= 4133) && (pixel_index <= 4153)) || ((pixel_index >= 4173) && (pixel_index <= 4176)) || ((pixel_index >= 4200) && (pixel_index <= 4217)) || ((pixel_index >= 4229) && (pixel_index <= 4251)) || ((pixel_index >= 4270) && (pixel_index <= 4272)) || ((pixel_index >= 4297) && (pixel_index <= 4313)) || ((pixel_index >= 4325) && (pixel_index <= 4347)) || ((pixel_index >= 4366) && (pixel_index <= 4367)) || ((pixel_index >= 4395) && (pixel_index <= 4408)) || ((pixel_index >= 4421) && (pixel_index <= 4453)) || pixel_index == 4492 || ((pixel_index >= 4499) && (pixel_index <= 4500)) || ((pixel_index >= 4517) && (pixel_index <= 4550)) || ((pixel_index >= 4613) && (pixel_index <= 4647)) || ((pixel_index >= 4674) && (pixel_index <= 4679)) || ((pixel_index >= 4709) && (pixel_index <= 4744)) || ((pixel_index >= 4769) && (pixel_index <= 4777)) || ((pixel_index >= 4805) && (pixel_index <= 4840)) || ((pixel_index >= 4864) && (pixel_index <= 4874)) || ((pixel_index >= 4901) && (pixel_index <= 4937)) || ((pixel_index >= 4960) && (pixel_index <= 4971)) || ((pixel_index >= 4997) && (pixel_index <= 5034)) || ((pixel_index >= 5055) && (pixel_index <= 5068)) || ((pixel_index >= 5093) && (pixel_index <= 5130)) || ((pixel_index >= 5151) && (pixel_index <= 5165)) || ((pixel_index >= 5189) && (pixel_index <= 5227)) || ((pixel_index >= 5247) && (pixel_index <= 5262)) || ((pixel_index >= 5285) && (pixel_index <= 5324)) || ((pixel_index >= 5343) && (pixel_index <= 5359)) || ((pixel_index >= 5381) && (pixel_index <= 5420)) || ((pixel_index >= 5438) && (pixel_index <= 5456)) || ((pixel_index >= 5477) && (pixel_index <= 5517)) || ((pixel_index >= 5534) && (pixel_index <= 5553)) || pixel_index == 5561 || ((pixel_index >= 5573) && (pixel_index <= 5614)) || ((pixel_index >= 5631) && (pixel_index <= 5650)) || ((pixel_index >= 5655) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5711)) || ((pixel_index >= 5727) && (pixel_index <= 5747)) || ((pixel_index >= 5750) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5807)) || ((pixel_index >= 5823) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5903)) || ((pixel_index >= 5920) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 5999)) || ((pixel_index >= 6017) && (pixel_index <= 6041)) || ((pixel_index >= 6053) && (pixel_index <= 6094)) || (pixel_index >= 6113) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 13) begin
            if (((pixel_index >= 5) && (pixel_index <= 69)) || ((pixel_index >= 80) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 163)) || ((pixel_index >= 177) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 258)) || ((pixel_index >= 273) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 350)) || ((pixel_index >= 369) && (pixel_index <= 377)) || ((pixel_index >= 389) && (pixel_index <= 443)) || ((pixel_index >= 465) && (pixel_index <= 473)) || ((pixel_index >= 485) && (pixel_index <= 537)) || ((pixel_index >= 561) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 632)) || ((pixel_index >= 656) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 727)) || ((pixel_index >= 750) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 822)) || ((pixel_index >= 847) && (pixel_index <= 857)) || ((pixel_index >= 869) && (pixel_index <= 918)) || ((pixel_index >= 947) && (pixel_index <= 953)) || ((pixel_index >= 965) && (pixel_index <= 1013)) || ((pixel_index >= 1044) && (pixel_index <= 1049)) || ((pixel_index >= 1061) && (pixel_index <= 1109)) || ((pixel_index >= 1138) && (pixel_index <= 1145)) || ((pixel_index >= 1157) && (pixel_index <= 1205)) || ((pixel_index >= 1233) && (pixel_index <= 1241)) || ((pixel_index >= 1253) && (pixel_index <= 1301)) || ((pixel_index >= 1329) && (pixel_index <= 1337)) || ((pixel_index >= 1349) && (pixel_index <= 1396)) || ((pixel_index >= 1425) && (pixel_index <= 1433)) || ((pixel_index >= 1445) && (pixel_index <= 1491)) || ((pixel_index >= 1521) && (pixel_index <= 1529)) || ((pixel_index >= 1541) && (pixel_index <= 1586)) || ((pixel_index >= 1617) && (pixel_index <= 1625)) || ((pixel_index >= 1637) && (pixel_index <= 1680)) || ((pixel_index >= 1712) && (pixel_index <= 1721)) || ((pixel_index >= 1733) && (pixel_index <= 1774)) || ((pixel_index >= 1808) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1870)) || ((pixel_index >= 1904) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 1967)) || ((pixel_index >= 2000) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2064)) || ((pixel_index >= 2097) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2163)) || ((pixel_index >= 2193) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2260)) || ((pixel_index >= 2290) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2360)) || ((pixel_index >= 2388) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2456)) || pixel_index == 2481 || ((pixel_index >= 2484) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2551)) || ((pixel_index >= 2577) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2648)) || ((pixel_index >= 2674) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2745)) || ((pixel_index >= 2768) && (pixel_index <= 2770)) || ((pixel_index >= 2772) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2841)) || ((pixel_index >= 2863) && (pixel_index <= 2866)) || ((pixel_index >= 2869) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2938)) || ((pixel_index >= 2957) && (pixel_index <= 2962)) || ((pixel_index >= 2966) && (pixel_index <= 2969)) || ((pixel_index >= 2981) && (pixel_index <= 3035)) || ((pixel_index >= 3053) && (pixel_index <= 3058)) || ((pixel_index >= 3063) && (pixel_index <= 3065)) || ((pixel_index >= 3077) && (pixel_index <= 3136)) || ((pixel_index >= 3147) && (pixel_index <= 3154)) || ((pixel_index >= 3160) && (pixel_index <= 3161)) || ((pixel_index >= 3173) && (pixel_index <= 3231)) || ((pixel_index >= 3240) && (pixel_index <= 3249)) || pixel_index == 3257 || ((pixel_index >= 3269) && (pixel_index <= 3327)) || ((pixel_index >= 3336) && (pixel_index <= 3345)) || ((pixel_index >= 3365) && (pixel_index <= 3421)) || ((pixel_index >= 3432) && (pixel_index <= 3441)) || ((pixel_index >= 3461) && (pixel_index <= 3516)) || ((pixel_index >= 3528) && (pixel_index <= 3537)) || ((pixel_index >= 3557) && (pixel_index <= 3579)) || ((pixel_index >= 3593) && (pixel_index <= 3611)) || ((pixel_index >= 3625) && (pixel_index <= 3632)) || ((pixel_index >= 3653) && (pixel_index <= 3675)) || ((pixel_index >= 3691) && (pixel_index <= 3705)) || ((pixel_index >= 3721) && (pixel_index <= 3728)) || ((pixel_index >= 3749) && (pixel_index <= 3771)) || ((pixel_index >= 3788) && (pixel_index <= 3799)) || ((pixel_index >= 3817) && (pixel_index <= 3823)) || ((pixel_index >= 3845) && (pixel_index <= 3868)) || ((pixel_index >= 3885) && (pixel_index <= 3895)) || ((pixel_index >= 3914) && (pixel_index <= 3919)) || ((pixel_index >= 3927) && (pixel_index <= 3928)) || ((pixel_index >= 3941) && (pixel_index <= 3965)) || ((pixel_index >= 3982) && (pixel_index <= 3991)) || ((pixel_index >= 4010) && (pixel_index <= 4014)) || ((pixel_index >= 4022) && (pixel_index <= 4025)) || ((pixel_index >= 4037) && (pixel_index <= 4062)) || ((pixel_index >= 4079) && (pixel_index <= 4086)) || ((pixel_index >= 4106) && (pixel_index <= 4109)) || ((pixel_index >= 4117) && (pixel_index <= 4121)) || ((pixel_index >= 4133) && (pixel_index <= 4158)) || ((pixel_index >= 4176) && (pixel_index <= 4181)) || ((pixel_index >= 4203) && (pixel_index <= 4204)) || ((pixel_index >= 4212) && (pixel_index <= 4217)) || ((pixel_index >= 4229) && (pixel_index <= 4256)) || ((pixel_index >= 4273) && (pixel_index <= 4277)) || ((pixel_index >= 4308) && (pixel_index <= 4313)) || ((pixel_index >= 4325) && (pixel_index <= 4353)) || ((pixel_index >= 4356) && (pixel_index <= 4359)) || ((pixel_index >= 4369) && (pixel_index <= 4372)) || ((pixel_index >= 4403) && (pixel_index <= 4409)) || ((pixel_index >= 4421) && (pixel_index <= 4455)) || ((pixel_index >= 4466) && (pixel_index <= 4467)) || ((pixel_index >= 4498) && (pixel_index <= 4505)) || ((pixel_index >= 4517) && (pixel_index <= 4552)) || ((pixel_index >= 4594) && (pixel_index <= 4601)) || ((pixel_index >= 4613) && (pixel_index <= 4649)) || ((pixel_index >= 4690) && (pixel_index <= 4697)) || ((pixel_index >= 4709) && (pixel_index <= 4745)) || pixel_index == 4786 || ((pixel_index >= 4788) && (pixel_index <= 4793)) || ((pixel_index >= 4805) && (pixel_index <= 4842)) || ((pixel_index >= 4887) && (pixel_index <= 4889)) || ((pixel_index >= 4901) && (pixel_index <= 4939)) || ((pixel_index >= 4966) && (pixel_index <= 4972)) || ((pixel_index >= 4997) && (pixel_index <= 5035)) || ((pixel_index >= 5061) && (pixel_index <= 5070)) || ((pixel_index >= 5093) && (pixel_index <= 5132)) || ((pixel_index >= 5157) && (pixel_index <= 5167)) || ((pixel_index >= 5189) && (pixel_index <= 5228)) || ((pixel_index >= 5253) && (pixel_index <= 5264)) || ((pixel_index >= 5285) && (pixel_index <= 5325)) || ((pixel_index >= 5348) && (pixel_index <= 5360)) || ((pixel_index >= 5381) && (pixel_index <= 5422)) || ((pixel_index >= 5444) && (pixel_index <= 5457)) || ((pixel_index >= 5477) && (pixel_index <= 5519)) || ((pixel_index >= 5540) && (pixel_index <= 5554)) || ((pixel_index >= 5573) && (pixel_index <= 5616)) || ((pixel_index >= 5636) && (pixel_index <= 5651)) || ((pixel_index >= 5669) && (pixel_index <= 5717)) || ((pixel_index >= 5732) && (pixel_index <= 5747)) || ((pixel_index >= 5765) && (pixel_index <= 5813)) || ((pixel_index >= 5828) && (pixel_index <= 5844)) || ((pixel_index >= 5861) && (pixel_index <= 5909)) || ((pixel_index >= 5924) && (pixel_index <= 5941)) || ((pixel_index >= 5957) && (pixel_index <= 6005)) || ((pixel_index >= 6020) && (pixel_index <= 6038)) || ((pixel_index >= 6053) && (pixel_index <= 6101)) || (pixel_index >= 6117) && (pixel_index <= 6134)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 14) begin
            if (((pixel_index >= 5) && (pixel_index <= 77)) || ((pixel_index >= 101) && (pixel_index <= 167)) || ((pixel_index >= 197) && (pixel_index <= 260)) || ((pixel_index >= 293) && (pixel_index <= 354)) || ((pixel_index >= 389) && (pixel_index <= 449)) || ((pixel_index >= 485) && (pixel_index <= 543)) || ((pixel_index >= 581) && (pixel_index <= 638)) || ((pixel_index >= 677) && (pixel_index <= 733)) || ((pixel_index >= 773) && (pixel_index <= 829)) || ((pixel_index >= 869) && (pixel_index <= 924)) || ((pixel_index >= 965) && (pixel_index <= 1020)) || ((pixel_index >= 1061) && (pixel_index <= 1116)) || ((pixel_index >= 1157) && (pixel_index <= 1211)) || ((pixel_index >= 1253) && (pixel_index <= 1307)) || ((pixel_index >= 1349) && (pixel_index <= 1401)) || ((pixel_index >= 1445) && (pixel_index <= 1495)) || ((pixel_index >= 1541) && (pixel_index <= 1588)) || ((pixel_index >= 1637) && (pixel_index <= 1683)) || ((pixel_index >= 1733) && (pixel_index <= 1779)) || ((pixel_index >= 1829) && (pixel_index <= 1876)) || ((pixel_index >= 1925) && (pixel_index <= 1973)) || ((pixel_index >= 2021) && (pixel_index <= 2070)) || ((pixel_index >= 2072) && (pixel_index <= 2073)) || ((pixel_index >= 2117) && (pixel_index <= 2169)) || ((pixel_index >= 2213) && (pixel_index <= 2265)) || ((pixel_index >= 2309) && (pixel_index <= 2362)) || ((pixel_index >= 2405) && (pixel_index <= 2461)) || ((pixel_index >= 2501) && (pixel_index <= 2558)) || ((pixel_index >= 2597) && (pixel_index <= 2653)) || ((pixel_index >= 2693) && (pixel_index <= 2749)) || ((pixel_index >= 2789) && (pixel_index <= 2846)) || ((pixel_index >= 2885) && (pixel_index <= 2942)) || ((pixel_index >= 2981) && (pixel_index <= 3039)) || ((pixel_index >= 3077) && (pixel_index <= 3136)) || ((pixel_index >= 3173) && (pixel_index <= 3232)) || pixel_index == 3257 || ((pixel_index >= 3269) && (pixel_index <= 3293)) || ((pixel_index >= 3300) && (pixel_index <= 3330)) || pixel_index == 3332 || ((pixel_index >= 3334) && (pixel_index <= 3335)) || pixel_index == 3350 || ((pixel_index >= 3352) && (pixel_index <= 3353)) || ((pixel_index >= 3365) && (pixel_index <= 3384)) || ((pixel_index >= 3400) && (pixel_index <= 3431)) || pixel_index == 3443 || ((pixel_index >= 3445) && (pixel_index <= 3449)) || ((pixel_index >= 3461) && (pixel_index <= 3480)) || ((pixel_index >= 3499) && (pixel_index <= 3526)) || ((pixel_index >= 3539) && (pixel_index <= 3545)) || ((pixel_index >= 3557) && (pixel_index <= 3576)) || ((pixel_index >= 3596) && (pixel_index <= 3622)) || pixel_index == 3632 || ((pixel_index >= 3634) && (pixel_index <= 3641)) || ((pixel_index >= 3653) && (pixel_index <= 3673)) || ((pixel_index >= 3693) && (pixel_index <= 3717)) || ((pixel_index >= 3728) && (pixel_index <= 3737)) || ((pixel_index >= 3749) && (pixel_index <= 3770)) || ((pixel_index >= 3790) && (pixel_index <= 3811)) || ((pixel_index >= 3824) && (pixel_index <= 3832)) || ((pixel_index >= 3845) && (pixel_index <= 3866)) || ((pixel_index >= 3886) && (pixel_index <= 3905)) || ((pixel_index >= 3921) && (pixel_index <= 3928)) || ((pixel_index >= 3941) && (pixel_index <= 3963)) || ((pixel_index >= 3983) && (pixel_index <= 3997)) || ((pixel_index >= 4017) && (pixel_index <= 4024)) || ((pixel_index >= 4037) && (pixel_index <= 4059)) || ((pixel_index >= 4080) && (pixel_index <= 4092)) || ((pixel_index >= 4114) && (pixel_index <= 4120)) || ((pixel_index >= 4133) && (pixel_index <= 4157)) || ((pixel_index >= 4177) && (pixel_index <= 4189)) || ((pixel_index >= 4210) && (pixel_index <= 4215)) || ((pixel_index >= 4229) && (pixel_index <= 4254)) || ((pixel_index >= 4257) && (pixel_index <= 4261)) || ((pixel_index >= 4274) && (pixel_index <= 4281)) || ((pixel_index >= 4306) && (pixel_index <= 4311)) || ((pixel_index >= 4325) && (pixel_index <= 4358)) || ((pixel_index >= 4370) && (pixel_index <= 4378)) || ((pixel_index >= 4402) && (pixel_index <= 4407)) || ((pixel_index >= 4421) && (pixel_index <= 4454)) || ((pixel_index >= 4467) && (pixel_index <= 4473)) || ((pixel_index >= 4499) && (pixel_index <= 4502)) || ((pixel_index >= 4517) && (pixel_index <= 4551)) || ((pixel_index >= 4564) && (pixel_index <= 4567)) || ((pixel_index >= 4594) && (pixel_index <= 4598)) || ((pixel_index >= 4613) && (pixel_index <= 4647)) || ((pixel_index >= 4660) && (pixel_index <= 4661)) || ((pixel_index >= 4691) && (pixel_index <= 4693)) || ((pixel_index >= 4709) && (pixel_index <= 4744)) || ((pixel_index >= 4805) && (pixel_index <= 4841)) || ((pixel_index >= 4901) && (pixel_index <= 4937)) || ((pixel_index >= 4997) && (pixel_index <= 5034)) || ((pixel_index >= 5093) && (pixel_index <= 5131)) || ((pixel_index >= 5189) && (pixel_index <= 5227)) || ((pixel_index >= 5285) && (pixel_index <= 5324)) || ((pixel_index >= 5381) && (pixel_index <= 5420)) || ((pixel_index >= 5477) && (pixel_index <= 5517)) || ((pixel_index >= 5573) && (pixel_index <= 5614)) || ((pixel_index >= 5646) && (pixel_index <= 5653)) || ((pixel_index >= 5669) && (pixel_index <= 5711)) || ((pixel_index >= 5722) && (pixel_index <= 5723)) || ((pixel_index >= 5742) && (pixel_index <= 5750)) || ((pixel_index >= 5765) && (pixel_index <= 5808)) || ((pixel_index >= 5815) && (pixel_index <= 5819)) || ((pixel_index >= 5837) && (pixel_index <= 5848)) || ((pixel_index >= 5861) && (pixel_index <= 5915)) || ((pixel_index >= 5933) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 6010)) || ((pixel_index >= 6029) && (pixel_index <= 6041)) || ((pixel_index >= 6053) && (pixel_index <= 6106)) || (pixel_index >= 6124) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 15) begin
            if (((pixel_index >= 5) && (pixel_index <= 82)) || ((pixel_index >= 101) && (pixel_index <= 177)) || ((pixel_index >= 197) && (pixel_index <= 264)) || ((pixel_index >= 293) && (pixel_index <= 357)) || ((pixel_index >= 389) && (pixel_index <= 451)) || ((pixel_index >= 485) && (pixel_index <= 546)) || ((pixel_index >= 581) && (pixel_index <= 641)) || ((pixel_index >= 677) && (pixel_index <= 736)) || ((pixel_index >= 773) && (pixel_index <= 831)) || ((pixel_index >= 869) && (pixel_index <= 926)) || ((pixel_index >= 965) && (pixel_index <= 1022)) || ((pixel_index >= 1061) && (pixel_index <= 1118)) || ((pixel_index >= 1157) && (pixel_index <= 1213)) || ((pixel_index >= 1253) && (pixel_index <= 1307)) || ((pixel_index >= 1349) && (pixel_index <= 1401)) || ((pixel_index >= 1445) && (pixel_index <= 1493)) || ((pixel_index >= 1541) && (pixel_index <= 1589)) || ((pixel_index >= 1637) && (pixel_index <= 1685)) || ((pixel_index >= 1733) && (pixel_index <= 1781)) || ((pixel_index >= 1829) && (pixel_index <= 1878)) || ((pixel_index >= 1925) && (pixel_index <= 1975)) || ((pixel_index >= 2021) && (pixel_index <= 2074)) || ((pixel_index >= 2117) && (pixel_index <= 2170)) || ((pixel_index >= 2213) && (pixel_index <= 2267)) || ((pixel_index >= 2309) && (pixel_index <= 2365)) || ((pixel_index >= 2405) && (pixel_index <= 2462)) || ((pixel_index >= 2501) && (pixel_index <= 2558)) || ((pixel_index >= 2597) && (pixel_index <= 2653)) || ((pixel_index >= 2693) && (pixel_index <= 2750)) || ((pixel_index >= 2789) && (pixel_index <= 2846)) || ((pixel_index >= 2885) && (pixel_index <= 2943)) || ((pixel_index >= 2981) && (pixel_index <= 3003)) || ((pixel_index >= 3005) && (pixel_index <= 3039)) || ((pixel_index >= 3077) && (pixel_index <= 3093)) || ((pixel_index >= 3107) && (pixel_index <= 3136)) || ((pixel_index >= 3173) && (pixel_index <= 3189)) || ((pixel_index >= 3206) && (pixel_index <= 3232)) || ((pixel_index >= 3269) && (pixel_index <= 3285)) || ((pixel_index >= 3305) && (pixel_index <= 3329)) || pixel_index == 3335 || ((pixel_index >= 3365) && (pixel_index <= 3382)) || ((pixel_index >= 3403) && (pixel_index <= 3431)) || ((pixel_index >= 3461) && (pixel_index <= 3479)) || ((pixel_index >= 3500) && (pixel_index <= 3527)) || pixel_index == 3543 || ((pixel_index >= 3557) && (pixel_index <= 3576)) || ((pixel_index >= 3596) && (pixel_index <= 3623)) || pixel_index == 3635 || ((pixel_index >= 3638) && (pixel_index <= 3641)) || ((pixel_index >= 3653) && (pixel_index <= 3672)) || ((pixel_index >= 3693) && (pixel_index <= 3718)) || ((pixel_index >= 3731) && (pixel_index <= 3732)) || ((pixel_index >= 3734) && (pixel_index <= 3737)) || ((pixel_index >= 3749) && (pixel_index <= 3769)) || ((pixel_index >= 3790) && (pixel_index <= 3814)) || ((pixel_index >= 3826) && (pixel_index <= 3832)) || ((pixel_index >= 3845) && (pixel_index <= 3865)) || ((pixel_index >= 3887) && (pixel_index <= 3909)) || ((pixel_index >= 3921) && (pixel_index <= 3928)) || ((pixel_index >= 3941) && (pixel_index <= 3963)) || ((pixel_index >= 3984) && (pixel_index <= 3997)) || ((pixel_index >= 4018) && (pixel_index <= 4024)) || ((pixel_index >= 4037) && (pixel_index <= 4064)) || ((pixel_index >= 4066) && (pixel_index <= 4067)) || ((pixel_index >= 4080) && (pixel_index <= 4093)) || ((pixel_index >= 4114) && (pixel_index <= 4120)) || ((pixel_index >= 4133) && (pixel_index <= 4164)) || ((pixel_index >= 4177) && (pixel_index <= 4186)) || ((pixel_index >= 4188) && (pixel_index <= 4189)) || ((pixel_index >= 4210) && (pixel_index <= 4216)) || ((pixel_index >= 4229) && (pixel_index <= 4260)) || ((pixel_index >= 4274) && (pixel_index <= 4282)) || ((pixel_index >= 4307) && (pixel_index <= 4311)) || ((pixel_index >= 4325) && (pixel_index <= 4357)) || ((pixel_index >= 4371) && (pixel_index <= 4377)) || ((pixel_index >= 4403) && (pixel_index <= 4407)) || ((pixel_index >= 4421) && (pixel_index <= 4454)) || ((pixel_index >= 4467) && (pixel_index <= 4470)) || ((pixel_index >= 4499) && (pixel_index <= 4503)) || ((pixel_index >= 4517) && (pixel_index <= 4550)) || pixel_index == 4564 || ((pixel_index >= 4595) && (pixel_index <= 4599)) || ((pixel_index >= 4613) && (pixel_index <= 4647)) || ((pixel_index >= 4691) && (pixel_index <= 4694)) || ((pixel_index >= 4709) && (pixel_index <= 4744)) || ((pixel_index >= 4787) && (pixel_index <= 4790)) || ((pixel_index >= 4805) && (pixel_index <= 4840)) || ((pixel_index >= 4884) && (pixel_index <= 4885)) || ((pixel_index >= 4901) && (pixel_index <= 4937)) || ((pixel_index >= 4997) && (pixel_index <= 5034)) || ((pixel_index >= 5093) && (pixel_index <= 5130)) || ((pixel_index >= 5189) && (pixel_index <= 5227)) || ((pixel_index >= 5285) && (pixel_index <= 5324)) || ((pixel_index >= 5381) && (pixel_index <= 5421)) || ((pixel_index >= 5477) && (pixel_index <= 5519)) || ((pixel_index >= 5529) && (pixel_index <= 5531)) || ((pixel_index >= 5573) && (pixel_index <= 5617)) || ((pixel_index >= 5619) && (pixel_index <= 5627)) || ((pixel_index >= 5669) && (pixel_index <= 5723)) || ((pixel_index >= 5743) && (pixel_index <= 5746)) || ((pixel_index >= 5765) && (pixel_index <= 5819)) || ((pixel_index >= 5838) && (pixel_index <= 5845)) || ((pixel_index >= 5861) && (pixel_index <= 5915)) || ((pixel_index >= 5934) && (pixel_index <= 5943)) || ((pixel_index >= 5957) && (pixel_index <= 6011)) || ((pixel_index >= 6030) && (pixel_index <= 6040)) || ((pixel_index >= 6053) && (pixel_index <= 6107)) || (pixel_index >= 6126) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 16) begin
            if (((pixel_index >= 5) && (pixel_index <= 87)) || ((pixel_index >= 101) && (pixel_index <= 181)) || ((pixel_index >= 197) && (pixel_index <= 267)) || ((pixel_index >= 293) && (pixel_index <= 360)) || ((pixel_index >= 389) && (pixel_index <= 453)) || ((pixel_index >= 485) && (pixel_index <= 548)) || ((pixel_index >= 581) && (pixel_index <= 642)) || ((pixel_index >= 677) && (pixel_index <= 738)) || ((pixel_index >= 773) && (pixel_index <= 833)) || ((pixel_index >= 869) && (pixel_index <= 928)) || ((pixel_index >= 965) && (pixel_index <= 1024)) || ((pixel_index >= 1061) && (pixel_index <= 1119)) || ((pixel_index >= 1157) && (pixel_index <= 1212)) || ((pixel_index >= 1253) && (pixel_index <= 1303)) || ((pixel_index >= 1349) && (pixel_index <= 1398)) || ((pixel_index >= 1445) && (pixel_index <= 1494)) || ((pixel_index >= 1541) && (pixel_index <= 1591)) || ((pixel_index >= 1637) && (pixel_index <= 1687)) || ((pixel_index >= 1733) && (pixel_index <= 1783)) || ((pixel_index >= 1829) && (pixel_index <= 1881)) || ((pixel_index >= 1925) && (pixel_index <= 1979)) || ((pixel_index >= 2021) && (pixel_index <= 2075)) || ((pixel_index >= 2117) && (pixel_index <= 2172)) || ((pixel_index >= 2213) && (pixel_index <= 2269)) || ((pixel_index >= 2309) && (pixel_index <= 2367)) || ((pixel_index >= 2405) && (pixel_index <= 2463)) || ((pixel_index >= 2501) && (pixel_index <= 2557)) || ((pixel_index >= 2597) && (pixel_index <= 2654)) || ((pixel_index >= 2693) && (pixel_index <= 2751)) || ((pixel_index >= 2789) && (pixel_index <= 2847)) || ((pixel_index >= 2885) && (pixel_index <= 2904)) || ((pixel_index >= 2913) && (pixel_index <= 2943)) || ((pixel_index >= 2981) && (pixel_index <= 2995)) || ((pixel_index >= 3011) && (pixel_index <= 3040)) || ((pixel_index >= 3077) && (pixel_index <= 3091)) || ((pixel_index >= 3110) && (pixel_index <= 3136)) || ((pixel_index >= 3173) && (pixel_index <= 3188)) || ((pixel_index >= 3209) && (pixel_index <= 3232)) || ((pixel_index >= 3269) && (pixel_index <= 3284)) || ((pixel_index >= 3306) && (pixel_index <= 3331)) || pixel_index == 3335 || ((pixel_index >= 3365) && (pixel_index <= 3381)) || ((pixel_index >= 3403) && (pixel_index <= 3431)) || ((pixel_index >= 3461) && (pixel_index <= 3478)) || ((pixel_index >= 3500) && (pixel_index <= 3527)) || ((pixel_index >= 3557) && (pixel_index <= 3575)) || ((pixel_index >= 3596) && (pixel_index <= 3623)) || ((pixel_index >= 3653) && (pixel_index <= 3671)) || ((pixel_index >= 3693) && (pixel_index <= 3719)) || pixel_index == 3731 || ((pixel_index >= 3734) && (pixel_index <= 3736)) || ((pixel_index >= 3749) && (pixel_index <= 3767)) || ((pixel_index >= 3790) && (pixel_index <= 3814)) || ((pixel_index >= 3827) && (pixel_index <= 3828)) || ((pixel_index >= 3830) && (pixel_index <= 3832)) || ((pixel_index >= 3845) && (pixel_index <= 3866)) || ((pixel_index >= 3887) && (pixel_index <= 3902)) || pixel_index == 3909 || ((pixel_index >= 3923) && (pixel_index <= 3928)) || ((pixel_index >= 3941) && (pixel_index <= 3964)) || pixel_index == 3970 || ((pixel_index >= 3984) && (pixel_index <= 3997)) || ((pixel_index >= 4018) && (pixel_index <= 4024)) || ((pixel_index >= 4037) && (pixel_index <= 4067)) || ((pixel_index >= 4081) && (pixel_index <= 4094)) || ((pixel_index >= 4114) && (pixel_index <= 4119)) || ((pixel_index >= 4133) && (pixel_index <= 4164)) || ((pixel_index >= 4178) && (pixel_index <= 4186)) || ((pixel_index >= 4210) && (pixel_index <= 4215)) || ((pixel_index >= 4229) && (pixel_index <= 4261)) || ((pixel_index >= 4274) && (pixel_index <= 4282)) || ((pixel_index >= 4307) && (pixel_index <= 4311)) || ((pixel_index >= 4325) && (pixel_index <= 4357)) || ((pixel_index >= 4371) && (pixel_index <= 4374)) || ((pixel_index >= 4403) && (pixel_index <= 4407)) || ((pixel_index >= 4421) && (pixel_index <= 4454)) || pixel_index == 4468 || ((pixel_index >= 4499) && (pixel_index <= 4503)) || ((pixel_index >= 4517) && (pixel_index <= 4551)) || ((pixel_index >= 4595) && (pixel_index <= 4598)) || ((pixel_index >= 4613) && (pixel_index <= 4648)) || ((pixel_index >= 4691) && (pixel_index <= 4694)) || ((pixel_index >= 4709) && (pixel_index <= 4744)) || ((pixel_index >= 4787) && (pixel_index <= 4790)) || ((pixel_index >= 4805) && (pixel_index <= 4841)) || ((pixel_index >= 4883) && (pixel_index <= 4886)) || ((pixel_index >= 4901) && (pixel_index <= 4938)) || pixel_index == 4981 || ((pixel_index >= 4997) && (pixel_index <= 5035)) || ((pixel_index >= 5093) && (pixel_index <= 5132)) || ((pixel_index >= 5189) && (pixel_index <= 5229)) || ((pixel_index >= 5285) && (pixel_index <= 5327)) || ((pixel_index >= 5338) && (pixel_index <= 5339)) || pixel_index == 5369 || ((pixel_index >= 5381) && (pixel_index <= 5435)) || ((pixel_index >= 5477) && (pixel_index <= 5531)) || ((pixel_index >= 5573) && (pixel_index <= 5627)) || ((pixel_index >= 5669) && (pixel_index <= 5723)) || pixel_index == 5743 || ((pixel_index >= 5765) && (pixel_index <= 5819)) || ((pixel_index >= 5839) && (pixel_index <= 5845)) || ((pixel_index >= 5861) && (pixel_index <= 5915)) || ((pixel_index >= 5934) && (pixel_index <= 5942)) || ((pixel_index >= 5957) && (pixel_index <= 6011)) || ((pixel_index >= 6030) && (pixel_index <= 6039)) || ((pixel_index >= 6053) && (pixel_index <= 6107)) || (pixel_index >= 6126) && (pixel_index <= 6136)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 17) begin
            if (((pixel_index >= 5) && (pixel_index <= 73)) || ((pixel_index >= 101) && (pixel_index <= 167)) || ((pixel_index >= 197) && (pixel_index <= 262)) || ((pixel_index >= 293) && (pixel_index <= 357)) || ((pixel_index >= 389) && (pixel_index <= 452)) || ((pixel_index >= 485) && (pixel_index <= 548)) || ((pixel_index >= 581) && (pixel_index <= 643)) || ((pixel_index >= 677) && (pixel_index <= 731)) || pixel_index == 735 || ((pixel_index >= 773) && (pixel_index <= 826)) || ((pixel_index >= 869) && (pixel_index <= 921)) || ((pixel_index >= 965) && (pixel_index <= 1017)) || ((pixel_index >= 1061) && (pixel_index <= 1114)) || ((pixel_index >= 1157) && (pixel_index <= 1210)) || ((pixel_index >= 1253) && (pixel_index <= 1306)) || ((pixel_index >= 1349) && (pixel_index <= 1402)) || ((pixel_index >= 1445) && (pixel_index <= 1501)) || ((pixel_index >= 1541) && (pixel_index <= 1598)) || ((pixel_index >= 1637) && (pixel_index <= 1694)) || ((pixel_index >= 1733) && (pixel_index <= 1791)) || ((pixel_index >= 1829) && (pixel_index <= 1889)) || ((pixel_index >= 1925) && (pixel_index <= 1985)) || ((pixel_index >= 2021) && (pixel_index <= 2081)) || ((pixel_index >= 2117) && (pixel_index <= 2176)) || ((pixel_index >= 2213) && (pixel_index <= 2272)) || ((pixel_index >= 2309) && (pixel_index <= 2369)) || ((pixel_index >= 2405) && (pixel_index <= 2465)) || ((pixel_index >= 2501) && (pixel_index <= 2561)) || ((pixel_index >= 2597) && (pixel_index <= 2614)) || ((pixel_index >= 2624) && (pixel_index <= 2658)) || ((pixel_index >= 2693) && (pixel_index <= 2710)) || ((pixel_index >= 2723) && (pixel_index <= 2754)) || ((pixel_index >= 2789) && (pixel_index <= 2804)) || ((pixel_index >= 2822) && (pixel_index <= 2850)) || ((pixel_index >= 2885) && (pixel_index <= 2899)) || ((pixel_index >= 2919) && (pixel_index <= 2949)) || ((pixel_index >= 2981) && (pixel_index <= 2995)) || ((pixel_index >= 3017) && (pixel_index <= 3049)) || ((pixel_index >= 3077) && (pixel_index <= 3091)) || ((pixel_index >= 3115) && (pixel_index <= 3145)) || ((pixel_index >= 3173) && (pixel_index <= 3188)) || ((pixel_index >= 3212) && (pixel_index <= 3241)) || ((pixel_index >= 3269) && (pixel_index <= 3285)) || ((pixel_index >= 3309) && (pixel_index <= 3337)) || ((pixel_index >= 3365) && (pixel_index <= 3382)) || ((pixel_index >= 3406) && (pixel_index <= 3433)) || pixel_index == 3449 || ((pixel_index >= 3461) && (pixel_index <= 3479)) || ((pixel_index >= 3503) && (pixel_index <= 3523)) || pixel_index == 3541 || ((pixel_index >= 3544) && (pixel_index <= 3545)) || ((pixel_index >= 3557) && (pixel_index <= 3574)) || ((pixel_index >= 3600) && (pixel_index <= 3616)) || ((pixel_index >= 3637) && (pixel_index <= 3641)) || ((pixel_index >= 3653) && (pixel_index <= 3674)) || ((pixel_index >= 3697) && (pixel_index <= 3712)) || ((pixel_index >= 3733) && (pixel_index <= 3737)) || ((pixel_index >= 3749) && (pixel_index <= 3771)) || ((pixel_index >= 3777) && (pixel_index <= 3779)) || ((pixel_index >= 3794) && (pixel_index <= 3804)) || ((pixel_index >= 3829) && (pixel_index <= 3833)) || ((pixel_index >= 3845) && (pixel_index <= 3876)) || ((pixel_index >= 3891) && (pixel_index <= 3900)) || ((pixel_index >= 3925) && (pixel_index <= 3929)) || ((pixel_index >= 3941) && (pixel_index <= 3973)) || ((pixel_index >= 3988) && (pixel_index <= 3994)) || ((pixel_index >= 4022) && (pixel_index <= 4025)) || ((pixel_index >= 4037) && (pixel_index <= 4070)) || ((pixel_index >= 4085) && (pixel_index <= 4087)) || ((pixel_index >= 4118) && (pixel_index <= 4121)) || ((pixel_index >= 4133) && (pixel_index <= 4167)) || ((pixel_index >= 4214) && (pixel_index <= 4217)) || ((pixel_index >= 4229) && (pixel_index <= 4264)) || ((pixel_index >= 4310) && (pixel_index <= 4313)) || ((pixel_index >= 4325) && (pixel_index <= 4361)) || ((pixel_index >= 4406) && (pixel_index <= 4409)) || ((pixel_index >= 4421) && (pixel_index <= 4458)) || ((pixel_index >= 4502) && (pixel_index <= 4505)) || ((pixel_index >= 4517) && (pixel_index <= 4555)) || ((pixel_index >= 4599) && (pixel_index <= 4601)) || ((pixel_index >= 4613) && (pixel_index <= 4652)) || ((pixel_index >= 4709) && (pixel_index <= 4749)) || ((pixel_index >= 4805) && (pixel_index <= 4847)) || ((pixel_index >= 4901) && (pixel_index <= 4945)) || ((pixel_index >= 4954) && (pixel_index <= 4957)) || ((pixel_index >= 4997) && (pixel_index <= 5053)) || ((pixel_index >= 5093) && (pixel_index <= 5149)) || ((pixel_index >= 5189) && (pixel_index <= 5245)) || ((pixel_index >= 5285) && (pixel_index <= 5341)) || ((pixel_index >= 5381) && (pixel_index <= 5437)) || ((pixel_index >= 5458) && (pixel_index <= 5463)) || ((pixel_index >= 5477) && (pixel_index <= 5533)) || ((pixel_index >= 5553) && (pixel_index <= 5560)) || ((pixel_index >= 5573) && (pixel_index <= 5629)) || ((pixel_index >= 5649) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5725)) || ((pixel_index >= 5745) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5821)) || ((pixel_index >= 5841) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5917)) || ((pixel_index >= 5936) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 6013)) || ((pixel_index >= 6032) && (pixel_index <= 6041)) || ((pixel_index >= 6053) && (pixel_index <= 6109)) || (pixel_index >= 6128) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 18) begin
            if (((pixel_index >= 5) && (pixel_index <= 81)) || ((pixel_index >= 101) && (pixel_index <= 177)) || ((pixel_index >= 197) && (pixel_index <= 274)) || ((pixel_index >= 293) && (pixel_index <= 371)) || ((pixel_index >= 389) && (pixel_index <= 468)) || ((pixel_index >= 485) && (pixel_index <= 564)) || ((pixel_index >= 581) && (pixel_index <= 660)) || ((pixel_index >= 677) && (pixel_index <= 756)) || ((pixel_index >= 773) && (pixel_index <= 853)) || ((pixel_index >= 869) && (pixel_index <= 949)) || ((pixel_index >= 965) && (pixel_index <= 1045)) || ((pixel_index >= 1061) && (pixel_index <= 1142)) || ((pixel_index >= 1157) && (pixel_index <= 1238)) || ((pixel_index >= 1253) && (pixel_index <= 1278)) || ((pixel_index >= 1283) && (pixel_index <= 1334)) || ((pixel_index >= 1349) && (pixel_index <= 1374)) || ((pixel_index >= 1381) && (pixel_index <= 1431)) || ((pixel_index >= 1445) && (pixel_index <= 1471)) || ((pixel_index >= 1480) && (pixel_index <= 1527)) || ((pixel_index >= 1541) && (pixel_index <= 1568)) || ((pixel_index >= 1579) && (pixel_index <= 1623)) || ((pixel_index >= 1637) && (pixel_index <= 1662)) || ((pixel_index >= 1678) && (pixel_index <= 1718)) || pixel_index == 1721 || ((pixel_index >= 1733) && (pixel_index <= 1750)) || ((pixel_index >= 1777) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1844)) || ((pixel_index >= 1875) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 1939)) || ((pixel_index >= 1972) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2036)) || ((pixel_index >= 2070) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2131)) || ((pixel_index >= 2167) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2227)) || ((pixel_index >= 2265) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2325)) || ((pixel_index >= 2362) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2421)) || ((pixel_index >= 2460) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2519)) || ((pixel_index >= 2558) && (pixel_index <= 2580)) || ((pixel_index >= 2597) && (pixel_index <= 2617)) || ((pixel_index >= 2655) && (pixel_index <= 2674)) || ((pixel_index >= 2693) && (pixel_index <= 2714)) || ((pixel_index >= 2753) && (pixel_index <= 2770)) || ((pixel_index >= 2789) && (pixel_index <= 2813)) || ((pixel_index >= 2850) && (pixel_index <= 2862)) || ((pixel_index >= 2864) && (pixel_index <= 2865)) || ((pixel_index >= 2885) && (pixel_index <= 2910)) || ((pixel_index >= 2947) && (pixel_index <= 2958)) || ((pixel_index >= 2981) && (pixel_index <= 3006)) || ((pixel_index >= 3022) && (pixel_index <= 3023)) || ((pixel_index >= 3045) && (pixel_index <= 3053)) || ((pixel_index >= 3077) && (pixel_index <= 3104)) || ((pixel_index >= 3116) && (pixel_index <= 3121)) || ((pixel_index >= 3142) && (pixel_index <= 3147)) || ((pixel_index >= 3173) && (pixel_index <= 3201)) || ((pixel_index >= 3210) && (pixel_index <= 3218)) || ((pixel_index >= 3239) && (pixel_index <= 3240)) || ((pixel_index >= 3269) && (pixel_index <= 3315)) || ((pixel_index >= 3365) && (pixel_index <= 3413)) || ((pixel_index >= 3461) && (pixel_index <= 3486)) || ((pixel_index >= 3498) && (pixel_index <= 3510)) || ((pixel_index >= 3557) && (pixel_index <= 3577)) || ((pixel_index >= 3595) && (pixel_index <= 3607)) || ((pixel_index >= 3653) && (pixel_index <= 3673)) || ((pixel_index >= 3691) && (pixel_index <= 3704)) || ((pixel_index >= 3749) && (pixel_index <= 3769)) || ((pixel_index >= 3786) && (pixel_index <= 3802)) || ((pixel_index >= 3845) && (pixel_index <= 3866)) || ((pixel_index >= 3882) && (pixel_index <= 3899)) || ((pixel_index >= 3941) && (pixel_index <= 3962)) || ((pixel_index >= 3977) && (pixel_index <= 3996)) || ((pixel_index >= 4037) && (pixel_index <= 4059)) || ((pixel_index >= 4072) && (pixel_index <= 4094)) || ((pixel_index >= 4133) && (pixel_index <= 4156)) || ((pixel_index >= 4167) && (pixel_index <= 4191)) || ((pixel_index >= 4229) && (pixel_index <= 4253)) || ((pixel_index >= 4263) && (pixel_index <= 4289)) || ((pixel_index >= 4325) && (pixel_index <= 4349)) || ((pixel_index >= 4359) && (pixel_index <= 4388)) || ((pixel_index >= 4396) && (pixel_index <= 4400)) || ((pixel_index >= 4421) && (pixel_index <= 4445)) || ((pixel_index >= 4455) && (pixel_index <= 4496)) || ((pixel_index >= 4517) && (pixel_index <= 4542)) || ((pixel_index >= 4550) && (pixel_index <= 4592)) || ((pixel_index >= 4613) && (pixel_index <= 4688)) || ((pixel_index >= 4709) && (pixel_index <= 4784)) || ((pixel_index >= 4805) && (pixel_index <= 4880)) || ((pixel_index >= 4901) && (pixel_index <= 4976)) || ((pixel_index >= 4997) && (pixel_index <= 5072)) || ((pixel_index >= 5093) && (pixel_index <= 5168)) || ((pixel_index >= 5189) && (pixel_index <= 5264)) || ((pixel_index >= 5285) && (pixel_index <= 5360)) || ((pixel_index >= 5381) && (pixel_index <= 5456)) || ((pixel_index >= 5477) && (pixel_index <= 5552)) || ((pixel_index >= 5573) && (pixel_index <= 5648)) || ((pixel_index >= 5669) && (pixel_index <= 5744)) || ((pixel_index >= 5765) && (pixel_index <= 5840)) || ((pixel_index >= 5861) && (pixel_index <= 5936)) || ((pixel_index >= 5957) && (pixel_index <= 6032)) || (pixel_index >= 6053) && (pixel_index <= 6128)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 19) begin
            if (((pixel_index >= 5) && (pixel_index <= 45)) || ((pixel_index >= 55) && (pixel_index <= 59)) || ((pixel_index >= 101) && (pixel_index <= 141)) || ((pixel_index >= 197) && (pixel_index <= 238)) || ((pixel_index >= 293) && (pixel_index <= 336)) || ((pixel_index >= 389) && (pixel_index <= 433)) || ((pixel_index >= 485) && (pixel_index <= 528)) || ((pixel_index >= 581) && (pixel_index <= 622)) || ((pixel_index >= 677) && (pixel_index <= 716)) || ((pixel_index >= 773) && (pixel_index <= 809)) || ((pixel_index >= 869) && (pixel_index <= 902)) || ((pixel_index >= 965) && (pixel_index <= 997)) || ((pixel_index >= 1061) && (pixel_index <= 1092)) || ((pixel_index >= 1157) && (pixel_index <= 1188)) || ((pixel_index >= 1253) && (pixel_index <= 1285)) || ((pixel_index >= 1304) && (pixel_index <= 1306)) || ((pixel_index >= 1349) && (pixel_index <= 1383)) || ((pixel_index >= 1398) && (pixel_index <= 1404)) || ((pixel_index >= 1445) && (pixel_index <= 1481)) || ((pixel_index >= 1492) && (pixel_index <= 1502)) || ((pixel_index >= 1541) && (pixel_index <= 1600)) || ((pixel_index >= 1637) && (pixel_index <= 1698)) || ((pixel_index >= 1733) && (pixel_index <= 1795)) || ((pixel_index >= 1829) && (pixel_index <= 1893)) || ((pixel_index >= 1925) && (pixel_index <= 1991)) || ((pixel_index >= 2021) && (pixel_index <= 2088)) || ((pixel_index >= 2117) && (pixel_index <= 2186)) || ((pixel_index >= 2213) && (pixel_index <= 2284)) || ((pixel_index >= 2309) && (pixel_index <= 2383)) || ((pixel_index >= 2405) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2969)) || ((pixel_index >= 2981) && (pixel_index <= 3065)) || ((pixel_index >= 3077) && (pixel_index <= 3161)) || ((pixel_index >= 3173) && (pixel_index <= 3257)) || ((pixel_index >= 3269) && (pixel_index <= 3353)) || ((pixel_index >= 3365) && (pixel_index <= 3449)) || ((pixel_index >= 3461) && (pixel_index <= 3545)) || ((pixel_index >= 3557) && (pixel_index <= 3641)) || ((pixel_index >= 3653) && (pixel_index <= 3737)) || ((pixel_index >= 3749) && (pixel_index <= 3833)) || ((pixel_index >= 3845) && (pixel_index <= 3929)) || ((pixel_index >= 3941) && (pixel_index <= 4025)) || ((pixel_index >= 4037) && (pixel_index <= 4121)) || ((pixel_index >= 4133) && (pixel_index <= 4217)) || ((pixel_index >= 4229) && (pixel_index <= 4313)) || ((pixel_index >= 4325) && (pixel_index <= 4409)) || ((pixel_index >= 4421) && (pixel_index <= 4505)) || ((pixel_index >= 4517) && (pixel_index <= 4601)) || ((pixel_index >= 4613) && (pixel_index <= 4697)) || ((pixel_index >= 4709) && (pixel_index <= 4793)) || ((pixel_index >= 4805) && (pixel_index <= 4889)) || ((pixel_index >= 4901) && (pixel_index <= 4985)) || ((pixel_index >= 4997) && (pixel_index <= 5081)) || ((pixel_index >= 5093) && (pixel_index <= 5177)) || ((pixel_index >= 5189) && (pixel_index <= 5215)) || ((pixel_index >= 5232) && (pixel_index <= 5273)) || ((pixel_index >= 5285) && (pixel_index <= 5308)) || ((pixel_index >= 5330) && (pixel_index <= 5369)) || ((pixel_index >= 5381) && (pixel_index <= 5403)) || ((pixel_index >= 5426) && (pixel_index <= 5465)) || ((pixel_index >= 5477) && (pixel_index <= 5498)) || ((pixel_index >= 5522) && (pixel_index <= 5561)) || ((pixel_index >= 5573) && (pixel_index <= 5595)) || ((pixel_index >= 5618) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5691)) || ((pixel_index >= 5714) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5787)) || ((pixel_index >= 5809) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5884)) || ((pixel_index >= 5905) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 5980)) || ((pixel_index >= 6000) && (pixel_index <= 6041)) || ((pixel_index >= 6053) && (pixel_index <= 6077)) || (pixel_index >= 6095) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 20) begin
            if (((pixel_index >= 5) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 377)) || ((pixel_index >= 389) && (pixel_index <= 473)) || ((pixel_index >= 485) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 857)) || ((pixel_index >= 869) && (pixel_index <= 953)) || ((pixel_index >= 965) && (pixel_index <= 1049)) || ((pixel_index >= 1061) && (pixel_index <= 1145)) || ((pixel_index >= 1157) && (pixel_index <= 1241)) || ((pixel_index >= 1253) && (pixel_index <= 1337)) || ((pixel_index >= 1349) && (pixel_index <= 1433)) || ((pixel_index >= 1445) && (pixel_index <= 1529)) || ((pixel_index >= 1541) && (pixel_index <= 1625)) || ((pixel_index >= 1637) && (pixel_index <= 1721)) || ((pixel_index >= 1733) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2969)) || ((pixel_index >= 2981) && (pixel_index <= 3065)) || ((pixel_index >= 3077) && (pixel_index <= 3161)) || ((pixel_index >= 3173) && (pixel_index <= 3257)) || ((pixel_index >= 3269) && (pixel_index <= 3353)) || ((pixel_index >= 3365) && (pixel_index <= 3449)) || ((pixel_index >= 3461) && (pixel_index <= 3545)) || ((pixel_index >= 3557) && (pixel_index <= 3641)) || ((pixel_index >= 3653) && (pixel_index <= 3737)) || ((pixel_index >= 3749) && (pixel_index <= 3833)) || ((pixel_index >= 3845) && (pixel_index <= 3929)) || ((pixel_index >= 3941) && (pixel_index <= 4025)) || ((pixel_index >= 4037) && (pixel_index <= 4121)) || ((pixel_index >= 4133) && (pixel_index <= 4217)) || ((pixel_index >= 4229) && (pixel_index <= 4313)) || ((pixel_index >= 4325) && (pixel_index <= 4409)) || ((pixel_index >= 4421) && (pixel_index <= 4505)) || ((pixel_index >= 4517) && (pixel_index <= 4601)) || ((pixel_index >= 4613) && (pixel_index <= 4653)) || ((pixel_index >= 4655) && (pixel_index <= 4656)) || pixel_index == 4659 || ((pixel_index >= 4661) && (pixel_index <= 4697)) || ((pixel_index >= 4709) && (pixel_index <= 4731)) || ((pixel_index >= 4759) && (pixel_index <= 4793)) || ((pixel_index >= 4805) && (pixel_index <= 4827)) || ((pixel_index >= 4855) && (pixel_index <= 4889)) || ((pixel_index >= 4901) && (pixel_index <= 4923)) || ((pixel_index >= 4950) && (pixel_index <= 4985)) || ((pixel_index >= 4997) && (pixel_index <= 5019)) || ((pixel_index >= 5046) && (pixel_index <= 5081)) || ((pixel_index >= 5093) && (pixel_index <= 5116)) || ((pixel_index >= 5142) && (pixel_index <= 5177)) || ((pixel_index >= 5189) && (pixel_index <= 5212)) || ((pixel_index >= 5238) && (pixel_index <= 5273)) || ((pixel_index >= 5285) && (pixel_index <= 5308)) || ((pixel_index >= 5333) && (pixel_index <= 5369)) || ((pixel_index >= 5381) && (pixel_index <= 5405)) || ((pixel_index >= 5428) && (pixel_index <= 5465)) || ((pixel_index >= 5477) && (pixel_index <= 5502)) || ((pixel_index >= 5523) && (pixel_index <= 5561)) || ((pixel_index >= 5573) && (pixel_index <= 5599)) || ((pixel_index >= 5618) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5696)) || ((pixel_index >= 5713) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5793)) || ((pixel_index >= 5809) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5889)) || ((pixel_index >= 5904) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 5986)) || ((pixel_index >= 6000) && (pixel_index <= 6041)) || ((pixel_index >= 6053) && (pixel_index <= 6082)) || (pixel_index >= 6096) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 21) begin
            if (((pixel_index >= 5) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 377)) || ((pixel_index >= 389) && (pixel_index <= 473)) || ((pixel_index >= 485) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 857)) || ((pixel_index >= 869) && (pixel_index <= 953)) || ((pixel_index >= 965) && (pixel_index <= 1049)) || ((pixel_index >= 1061) && (pixel_index <= 1145)) || ((pixel_index >= 1157) && (pixel_index <= 1241)) || ((pixel_index >= 1253) && (pixel_index <= 1337)) || ((pixel_index >= 1349) && (pixel_index <= 1433)) || ((pixel_index >= 1445) && (pixel_index <= 1529)) || ((pixel_index >= 1541) && (pixel_index <= 1625)) || ((pixel_index >= 1637) && (pixel_index <= 1721)) || ((pixel_index >= 1733) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2149)) || ((pixel_index >= 2164) && (pixel_index <= 2168)) || ((pixel_index >= 2171) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2242)) || pixel_index == 2263 || ((pixel_index >= 2268) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2337)) || pixel_index == 2362 || ((pixel_index >= 2365) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2432)) || ((pixel_index >= 2460) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2528)) || ((pixel_index >= 2556) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2624)) || ((pixel_index >= 2652) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2720)) || ((pixel_index >= 2748) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2817)) || ((pixel_index >= 2843) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2913)) || ((pixel_index >= 2939) && (pixel_index <= 2969)) || ((pixel_index >= 2981) && (pixel_index <= 3009)) || ((pixel_index >= 3034) && (pixel_index <= 3065)) || ((pixel_index >= 3077) && (pixel_index <= 3106)) || ((pixel_index >= 3130) && (pixel_index <= 3161)) || ((pixel_index >= 3173) && (pixel_index <= 3202)) || ((pixel_index >= 3225) && (pixel_index <= 3257)) || ((pixel_index >= 3269) && (pixel_index <= 3299)) || ((pixel_index >= 3320) && (pixel_index <= 3353)) || ((pixel_index >= 3365) && (pixel_index <= 3396)) || ((pixel_index >= 3415) && (pixel_index <= 3449)) || ((pixel_index >= 3461) && (pixel_index <= 3493)) || ((pixel_index >= 3510) && (pixel_index <= 3545)) || ((pixel_index >= 3557) && (pixel_index <= 3590)) || ((pixel_index >= 3605) && (pixel_index <= 3641)) || ((pixel_index >= 3653) && (pixel_index <= 3686)) || ((pixel_index >= 3701) && (pixel_index <= 3737)) || ((pixel_index >= 3749) && (pixel_index <= 3782)) || ((pixel_index >= 3796) && (pixel_index <= 3833)) || ((pixel_index >= 3845) && (pixel_index <= 3878)) || ((pixel_index >= 3892) && (pixel_index <= 3929)) || ((pixel_index >= 3941) && (pixel_index <= 3974)) || ((pixel_index >= 3988) && (pixel_index <= 4025)) || ((pixel_index >= 4037) && (pixel_index <= 4070)) || ((pixel_index >= 4084) && (pixel_index <= 4121)) || ((pixel_index >= 4133) && (pixel_index <= 4168)) || ((pixel_index >= 4179) && (pixel_index <= 4217)) || ((pixel_index >= 4229) && (pixel_index <= 4313)) || ((pixel_index >= 4325) && (pixel_index <= 4409)) || ((pixel_index >= 4421) && (pixel_index <= 4505)) || ((pixel_index >= 4517) && (pixel_index <= 4601)) || ((pixel_index >= 4613) && (pixel_index <= 4697)) || ((pixel_index >= 4709) && (pixel_index <= 4793)) || ((pixel_index >= 4805) && (pixel_index <= 4889)) || ((pixel_index >= 4901) && (pixel_index <= 4985)) || ((pixel_index >= 4997) && (pixel_index <= 5081)) || ((pixel_index >= 5093) && (pixel_index <= 5177)) || ((pixel_index >= 5189) && (pixel_index <= 5273)) || ((pixel_index >= 5285) && (pixel_index <= 5369)) || ((pixel_index >= 5381) && (pixel_index <= 5465)) || ((pixel_index >= 5477) && (pixel_index <= 5561)) || ((pixel_index >= 5573) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 6041)) || (pixel_index >= 6053) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 22) begin
            if (((pixel_index >= 5) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 377)) || ((pixel_index >= 389) && (pixel_index <= 473)) || ((pixel_index >= 485) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 614)) || ((pixel_index >= 627) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 707)) || ((pixel_index >= 726) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 802)) || ((pixel_index >= 824) && (pixel_index <= 857)) || ((pixel_index >= 869) && (pixel_index <= 898)) || ((pixel_index >= 922) && (pixel_index <= 924)) || ((pixel_index >= 927) && (pixel_index <= 953)) || ((pixel_index >= 965) && (pixel_index <= 994)) || ((pixel_index >= 1024) && (pixel_index <= 1049)) || ((pixel_index >= 1061) && (pixel_index <= 1090)) || ((pixel_index >= 1116) && (pixel_index <= 1118)) || ((pixel_index >= 1120) && (pixel_index <= 1145)) || ((pixel_index >= 1157) && (pixel_index <= 1186)) || ((pixel_index >= 1212) && (pixel_index <= 1214)) || ((pixel_index >= 1216) && (pixel_index <= 1241)) || ((pixel_index >= 1253) && (pixel_index <= 1282)) || ((pixel_index >= 1308) && (pixel_index <= 1310)) || ((pixel_index >= 1312) && (pixel_index <= 1337)) || ((pixel_index >= 1349) && (pixel_index <= 1378)) || ((pixel_index >= 1404) && (pixel_index <= 1405)) || ((pixel_index >= 1407) && (pixel_index <= 1433)) || ((pixel_index >= 1445) && (pixel_index <= 1474)) || pixel_index == 1500 || ((pixel_index >= 1503) && (pixel_index <= 1529)) || ((pixel_index >= 1541) && (pixel_index <= 1571)) || ((pixel_index >= 1598) && (pixel_index <= 1625)) || ((pixel_index >= 1637) && (pixel_index <= 1667)) || ((pixel_index >= 1692) && (pixel_index <= 1721)) || ((pixel_index >= 1733) && (pixel_index <= 1764)) || ((pixel_index >= 1787) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1861)) || ((pixel_index >= 1881) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 1958)) || ((pixel_index >= 1976) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2054)) || ((pixel_index >= 2071) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2151)) || ((pixel_index >= 2165) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2247)) || ((pixel_index >= 2261) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2342)) || ((pixel_index >= 2356) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2438)) || ((pixel_index >= 2452) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2535)) || ((pixel_index >= 2548) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2632)) || ((pixel_index >= 2644) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2733)) || ((pixel_index >= 2738) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2969)) || ((pixel_index >= 2981) && (pixel_index <= 3065)) || ((pixel_index >= 3077) && (pixel_index <= 3161)) || ((pixel_index >= 3173) && (pixel_index <= 3257)) || ((pixel_index >= 3269) && (pixel_index <= 3353)) || ((pixel_index >= 3365) && (pixel_index <= 3449)) || ((pixel_index >= 3461) && (pixel_index <= 3545)) || ((pixel_index >= 3557) && (pixel_index <= 3641)) || ((pixel_index >= 3653) && (pixel_index <= 3737)) || ((pixel_index >= 3749) && (pixel_index <= 3833)) || ((pixel_index >= 3845) && (pixel_index <= 3929)) || ((pixel_index >= 3941) && (pixel_index <= 4025)) || ((pixel_index >= 4037) && (pixel_index <= 4121)) || ((pixel_index >= 4133) && (pixel_index <= 4217)) || ((pixel_index >= 4229) && (pixel_index <= 4313)) || ((pixel_index >= 4325) && (pixel_index <= 4409)) || ((pixel_index >= 4421) && (pixel_index <= 4505)) || ((pixel_index >= 4517) && (pixel_index <= 4601)) || ((pixel_index >= 4613) && (pixel_index <= 4697)) || ((pixel_index >= 4709) && (pixel_index <= 4793)) || ((pixel_index >= 4805) && (pixel_index <= 4889)) || ((pixel_index >= 4901) && (pixel_index <= 4985)) || ((pixel_index >= 4997) && (pixel_index <= 5081)) || ((pixel_index >= 5093) && (pixel_index <= 5177)) || ((pixel_index >= 5189) && (pixel_index <= 5273)) || ((pixel_index >= 5285) && (pixel_index <= 5369)) || ((pixel_index >= 5381) && (pixel_index <= 5465)) || ((pixel_index >= 5477) && (pixel_index <= 5561)) || ((pixel_index >= 5573) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 6041)) || (pixel_index >= 6053) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 23) begin
            if (((pixel_index >= 5) && (pixel_index <= 34)) || ((pixel_index >= 49) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 130)) || ((pixel_index >= 148) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 226)) || ((pixel_index >= 247) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 321)) || ((pixel_index >= 345) && (pixel_index <= 377)) || ((pixel_index >= 389) && (pixel_index <= 417)) || ((pixel_index >= 443) && (pixel_index <= 473)) || ((pixel_index >= 485) && (pixel_index <= 514)) || ((pixel_index >= 540) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 610)) || ((pixel_index >= 640) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 706)) || ((pixel_index >= 734) && (pixel_index <= 735)) || ((pixel_index >= 737) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 802)) || ((pixel_index >= 829) && (pixel_index <= 832)) || ((pixel_index >= 834) && (pixel_index <= 857)) || ((pixel_index >= 869) && (pixel_index <= 899)) || ((pixel_index >= 925) && (pixel_index <= 928)) || ((pixel_index >= 930) && (pixel_index <= 953)) || ((pixel_index >= 965) && (pixel_index <= 995)) || ((pixel_index >= 1020) && (pixel_index <= 1023)) || ((pixel_index >= 1025) && (pixel_index <= 1049)) || ((pixel_index >= 1061) && (pixel_index <= 1092)) || ((pixel_index >= 1115) && (pixel_index <= 1118)) || ((pixel_index >= 1121) && (pixel_index <= 1145)) || ((pixel_index >= 1157) && (pixel_index <= 1189)) || ((pixel_index >= 1210) && (pixel_index <= 1213)) || ((pixel_index >= 1216) && (pixel_index <= 1241)) || ((pixel_index >= 1253) && (pixel_index <= 1285)) || ((pixel_index >= 1306) && (pixel_index <= 1307)) || ((pixel_index >= 1311) && (pixel_index <= 1337)) || ((pixel_index >= 1349) && (pixel_index <= 1382)) || ((pixel_index >= 1404) && (pixel_index <= 1433)) || ((pixel_index >= 1445) && (pixel_index <= 1478)) || ((pixel_index >= 1495) && (pixel_index <= 1529)) || ((pixel_index >= 1541) && (pixel_index <= 1574)) || ((pixel_index >= 1590) && (pixel_index <= 1625)) || ((pixel_index >= 1637) && (pixel_index <= 1669)) || ((pixel_index >= 1684) && (pixel_index <= 1721)) || ((pixel_index >= 1733) && (pixel_index <= 1765)) || ((pixel_index >= 1779) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1861)) || ((pixel_index >= 1875) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 1959)) || ((pixel_index >= 1971) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2058)) || ((pixel_index >= 2067) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2969)) || ((pixel_index >= 2981) && (pixel_index <= 3065)) || ((pixel_index >= 3077) && (pixel_index <= 3161)) || ((pixel_index >= 3173) && (pixel_index <= 3257)) || ((pixel_index >= 3269) && (pixel_index <= 3353)) || ((pixel_index >= 3365) && (pixel_index <= 3449)) || ((pixel_index >= 3461) && (pixel_index <= 3545)) || ((pixel_index >= 3557) && (pixel_index <= 3641)) || ((pixel_index >= 3653) && (pixel_index <= 3737)) || ((pixel_index >= 3749) && (pixel_index <= 3833)) || ((pixel_index >= 3845) && (pixel_index <= 3929)) || ((pixel_index >= 3941) && (pixel_index <= 4025)) || ((pixel_index >= 4037) && (pixel_index <= 4121)) || ((pixel_index >= 4133) && (pixel_index <= 4217)) || ((pixel_index >= 4229) && (pixel_index <= 4313)) || ((pixel_index >= 4325) && (pixel_index <= 4409)) || ((pixel_index >= 4421) && (pixel_index <= 4505)) || ((pixel_index >= 4517) && (pixel_index <= 4601)) || ((pixel_index >= 4613) && (pixel_index <= 4697)) || ((pixel_index >= 4709) && (pixel_index <= 4793)) || ((pixel_index >= 4805) && (pixel_index <= 4889)) || ((pixel_index >= 4901) && (pixel_index <= 4985)) || ((pixel_index >= 4997) && (pixel_index <= 5081)) || ((pixel_index >= 5093) && (pixel_index <= 5177)) || ((pixel_index >= 5189) && (pixel_index <= 5273)) || ((pixel_index >= 5285) && (pixel_index <= 5369)) || ((pixel_index >= 5381) && (pixel_index <= 5465)) || ((pixel_index >= 5477) && (pixel_index <= 5561)) || ((pixel_index >= 5573) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 6041)) || (pixel_index >= 6053) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 24) begin
            if (((pixel_index >= 5) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 377)) || ((pixel_index >= 389) && (pixel_index <= 473)) || ((pixel_index >= 485) && (pixel_index <= 515)) || ((pixel_index >= 519) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 610)) || ((pixel_index >= 620) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 705)) || ((pixel_index >= 720) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 801)) || ((pixel_index >= 819) && (pixel_index <= 857)) || ((pixel_index >= 869) && (pixel_index <= 897)) || ((pixel_index >= 918) && (pixel_index <= 953)) || ((pixel_index >= 965) && (pixel_index <= 993)) || ((pixel_index >= 1016) && (pixel_index <= 1049)) || ((pixel_index >= 1061) && (pixel_index <= 1089)) || ((pixel_index >= 1115) && (pixel_index <= 1145)) || ((pixel_index >= 1157) && (pixel_index <= 1185)) || ((pixel_index >= 1212) && (pixel_index <= 1241)) || ((pixel_index >= 1253) && (pixel_index <= 1282)) || ((pixel_index >= 1309) && (pixel_index <= 1337)) || ((pixel_index >= 1349) && (pixel_index <= 1378)) || ((pixel_index >= 1410) && (pixel_index <= 1433)) || ((pixel_index >= 1445) && (pixel_index <= 1475)) || ((pixel_index >= 1506) && (pixel_index <= 1529)) || ((pixel_index >= 1541) && (pixel_index <= 1571)) || ((pixel_index >= 1598) && (pixel_index <= 1600)) || ((pixel_index >= 1603) && (pixel_index <= 1625)) || ((pixel_index >= 1637) && (pixel_index <= 1668)) || ((pixel_index >= 1694) && (pixel_index <= 1697)) || ((pixel_index >= 1699) && (pixel_index <= 1721)) || ((pixel_index >= 1733) && (pixel_index <= 1765)) || pixel_index == 1788 || ((pixel_index >= 1790) && (pixel_index <= 1792)) || ((pixel_index >= 1795) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1861)) || ((pixel_index >= 1883) && (pixel_index <= 1888)) || ((pixel_index >= 1890) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 1957)) || ((pixel_index >= 1978) && (pixel_index <= 1982)) || ((pixel_index >= 1986) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2053)) || ((pixel_index >= 2074) && (pixel_index <= 2075)) || ((pixel_index >= 2081) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2149)) || ((pixel_index >= 2175) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2244)) || ((pixel_index >= 2264) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2340)) || ((pixel_index >= 2357) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2436)) || ((pixel_index >= 2451) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2534)) || ((pixel_index >= 2547) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2633)) || ((pixel_index >= 2643) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2733)) || ((pixel_index >= 2738) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2969)) || ((pixel_index >= 2981) && (pixel_index <= 3065)) || ((pixel_index >= 3077) && (pixel_index <= 3161)) || ((pixel_index >= 3173) && (pixel_index <= 3257)) || ((pixel_index >= 3269) && (pixel_index <= 3353)) || ((pixel_index >= 3365) && (pixel_index <= 3449)) || ((pixel_index >= 3461) && (pixel_index <= 3545)) || ((pixel_index >= 3557) && (pixel_index <= 3641)) || ((pixel_index >= 3653) && (pixel_index <= 3737)) || ((pixel_index >= 3749) && (pixel_index <= 3833)) || ((pixel_index >= 3845) && (pixel_index <= 3929)) || ((pixel_index >= 3941) && (pixel_index <= 4025)) || ((pixel_index >= 4037) && (pixel_index <= 4121)) || ((pixel_index >= 4133) && (pixel_index <= 4217)) || ((pixel_index >= 4229) && (pixel_index <= 4313)) || ((pixel_index >= 4325) && (pixel_index <= 4409)) || ((pixel_index >= 4421) && (pixel_index <= 4505)) || ((pixel_index >= 4517) && (pixel_index <= 4601)) || ((pixel_index >= 4613) && (pixel_index <= 4697)) || ((pixel_index >= 4709) && (pixel_index <= 4793)) || ((pixel_index >= 4805) && (pixel_index <= 4889)) || ((pixel_index >= 4901) && (pixel_index <= 4985)) || ((pixel_index >= 4997) && (pixel_index <= 5081)) || ((pixel_index >= 5093) && (pixel_index <= 5177)) || ((pixel_index >= 5189) && (pixel_index <= 5273)) || ((pixel_index >= 5285) && (pixel_index <= 5369)) || ((pixel_index >= 5381) && (pixel_index <= 5465)) || ((pixel_index >= 5477) && (pixel_index <= 5561)) || ((pixel_index >= 5573) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 6041)) || (pixel_index >= 6053) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 25) begin
            if (((pixel_index >= 5) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 377)) || ((pixel_index >= 389) && (pixel_index <= 473)) || ((pixel_index >= 485) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 857)) || ((pixel_index >= 869) && (pixel_index <= 953)) || ((pixel_index >= 965) && (pixel_index <= 1049)) || ((pixel_index >= 1061) && (pixel_index <= 1145)) || ((pixel_index >= 1157) && (pixel_index <= 1241)) || ((pixel_index >= 1253) && (pixel_index <= 1337)) || ((pixel_index >= 1349) && (pixel_index <= 1433)) || ((pixel_index >= 1445) && (pixel_index <= 1529)) || ((pixel_index >= 1541) && (pixel_index <= 1625)) || ((pixel_index >= 1637) && (pixel_index <= 1721)) || ((pixel_index >= 1733) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2818)) || ((pixel_index >= 2823) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2913)) || ((pixel_index >= 2923) && (pixel_index <= 2969)) || ((pixel_index >= 2981) && (pixel_index <= 3009)) || ((pixel_index >= 3023) && (pixel_index <= 3065)) || ((pixel_index >= 3077) && (pixel_index <= 3105)) || ((pixel_index >= 3122) && (pixel_index <= 3161)) || ((pixel_index >= 3173) && (pixel_index <= 3201)) || ((pixel_index >= 3220) && (pixel_index <= 3257)) || ((pixel_index >= 3269) && (pixel_index <= 3297)) || ((pixel_index >= 3319) && (pixel_index <= 3353)) || ((pixel_index >= 3365) && (pixel_index <= 3393)) || ((pixel_index >= 3417) && (pixel_index <= 3449)) || ((pixel_index >= 3461) && (pixel_index <= 3489)) || ((pixel_index >= 3515) && (pixel_index <= 3545)) || ((pixel_index >= 3557) && (pixel_index <= 3585)) || ((pixel_index >= 3613) && (pixel_index <= 3641)) || ((pixel_index >= 3653) && (pixel_index <= 3682)) || ((pixel_index >= 3710) && (pixel_index <= 3737)) || ((pixel_index >= 3749) && (pixel_index <= 3778)) || ((pixel_index >= 3810) && (pixel_index <= 3833)) || ((pixel_index >= 3845) && (pixel_index <= 3875)) || ((pixel_index >= 3907) && (pixel_index <= 3929)) || ((pixel_index >= 3941) && (pixel_index <= 3972)) || ((pixel_index >= 3999) && (pixel_index <= 4001)) || ((pixel_index >= 4003) && (pixel_index <= 4025)) || ((pixel_index >= 4037) && (pixel_index <= 4068)) || ((pixel_index >= 4094) && (pixel_index <= 4097)) || ((pixel_index >= 4099) && (pixel_index <= 4121)) || ((pixel_index >= 4133) && (pixel_index <= 4164)) || ((pixel_index >= 4189) && (pixel_index <= 4192)) || ((pixel_index >= 4195) && (pixel_index <= 4217)) || ((pixel_index >= 4229) && (pixel_index <= 4260)) || ((pixel_index >= 4284) && (pixel_index <= 4288)) || ((pixel_index >= 4291) && (pixel_index <= 4313)) || ((pixel_index >= 4325) && (pixel_index <= 4356)) || ((pixel_index >= 4379) && (pixel_index <= 4382)) || ((pixel_index >= 4386) && (pixel_index <= 4409)) || ((pixel_index >= 4421) && (pixel_index <= 4452)) || ((pixel_index >= 4474) && (pixel_index <= 4475)) || ((pixel_index >= 4481) && (pixel_index <= 4505)) || ((pixel_index >= 4517) && (pixel_index <= 4548)) || ((pixel_index >= 4575) && (pixel_index <= 4601)) || ((pixel_index >= 4613) && (pixel_index <= 4644)) || ((pixel_index >= 4662) && (pixel_index <= 4697)) || ((pixel_index >= 4709) && (pixel_index <= 4740)) || ((pixel_index >= 4755) && (pixel_index <= 4793)) || ((pixel_index >= 4805) && (pixel_index <= 4836)) || ((pixel_index >= 4851) && (pixel_index <= 4889)) || ((pixel_index >= 4901) && (pixel_index <= 4933)) || ((pixel_index >= 4946) && (pixel_index <= 4985)) || ((pixel_index >= 4997) && (pixel_index <= 5031)) || ((pixel_index >= 5042) && (pixel_index <= 5081)) || ((pixel_index >= 5093) && (pixel_index <= 5130)) || ((pixel_index >= 5138) && (pixel_index <= 5177)) || ((pixel_index >= 5189) && (pixel_index <= 5273)) || ((pixel_index >= 5285) && (pixel_index <= 5369)) || ((pixel_index >= 5381) && (pixel_index <= 5465)) || ((pixel_index >= 5477) && (pixel_index <= 5561)) || ((pixel_index >= 5573) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 6041)) || (pixel_index >= 6053) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 26) begin
            if (((pixel_index >= 3678) && (pixel_index <= 3689)) || ((pixel_index >= 3774) && (pixel_index <= 3785)) || ((pixel_index >= 3791) && (pixel_index <= 3793)) || ((pixel_index >= 3870) && (pixel_index <= 3881)) || ((pixel_index >= 3887) && (pixel_index <= 3891)) || ((pixel_index >= 3966) && (pixel_index <= 3978)) || ((pixel_index >= 3983) && (pixel_index <= 3989)) || ((pixel_index >= 4062) && (pixel_index <= 4074)) || ((pixel_index >= 4078) && (pixel_index <= 4088)) || ((pixel_index >= 4158) && (pixel_index <= 4170)) || ((pixel_index >= 4174) && (pixel_index <= 4186)) || ((pixel_index >= 4254) && (pixel_index <= 4267)) || ((pixel_index >= 4270) && (pixel_index <= 4282)) || ((pixel_index >= 4351) && (pixel_index <= 4363)) || ((pixel_index >= 4366) && (pixel_index <= 4378)) || pixel_index == 4380 || ((pixel_index >= 4447) && (pixel_index <= 4460)) || ((pixel_index >= 4463) && (pixel_index <= 4474)) || ((pixel_index >= 4476) && (pixel_index <= 4478)) || ((pixel_index >= 4543) && (pixel_index <= 4548)) || ((pixel_index >= 4550) && (pixel_index <= 4557)) || ((pixel_index >= 4559) && (pixel_index <= 4569)) || ((pixel_index >= 4571) && (pixel_index <= 4575)) || ((pixel_index >= 4640) && (pixel_index <= 4645)) || ((pixel_index >= 4647) && (pixel_index <= 4665)) || ((pixel_index >= 4667) && (pixel_index <= 4672)) || ((pixel_index >= 4736) && (pixel_index <= 4742)) || ((pixel_index >= 4744) && (pixel_index <= 4760)) || ((pixel_index >= 4762) && (pixel_index <= 4770)) || ((pixel_index >= 4833) && (pixel_index <= 4853)) || ((pixel_index >= 4858) && (pixel_index <= 4867)) || ((pixel_index >= 4930) && (pixel_index <= 4951)) || ((pixel_index >= 4953) && (pixel_index <= 4965)) || ((pixel_index >= 5027) && (pixel_index <= 5063)) || ((pixel_index >= 5123) && (pixel_index <= 5156)) || ((pixel_index >= 5158) && (pixel_index <= 5160)) || ((pixel_index >= 5220) && (pixel_index <= 5251)) || ((pixel_index >= 5255) && (pixel_index <= 5256)) || ((pixel_index >= 5316) && (pixel_index <= 5347)) || ((pixel_index >= 5351) && (pixel_index <= 5352)) || ((pixel_index >= 5412) && (pixel_index <= 5441)) || ((pixel_index >= 5446) && (pixel_index <= 5448)) || ((pixel_index >= 5507) && (pixel_index <= 5536)) || ((pixel_index >= 5540) && (pixel_index <= 5543)) || ((pixel_index >= 5602) && (pixel_index <= 5638)) || ((pixel_index >= 5698) && (pixel_index <= 5721)) || ((pixel_index >= 5723) && (pixel_index <= 5733)) || ((pixel_index >= 5795) && (pixel_index <= 5815)) || ((pixel_index >= 5891) && (pixel_index <= 5909)) || ((pixel_index >= 5988) && (pixel_index <= 6004)) || (pixel_index >= 6085) && (pixel_index <= 6099)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 27) begin
            if (((pixel_index >= 3015) && (pixel_index <= 3017)) || ((pixel_index >= 3111) && (pixel_index <= 3113)) || ((pixel_index >= 3206) && (pixel_index <= 3208)) || ((pixel_index >= 3301) && (pixel_index <= 3303)) || ((pixel_index >= 3396) && (pixel_index <= 3398)) || ((pixel_index >= 3491) && (pixel_index <= 3493)) || pixel_index == 3580 || ((pixel_index >= 3584) && (pixel_index <= 3588)) || ((pixel_index >= 3602) && (pixel_index <= 3603)) || ((pixel_index >= 3675) && (pixel_index <= 3676)) || ((pixel_index >= 3679) && (pixel_index <= 3683)) || ((pixel_index >= 3697) && (pixel_index <= 3701)) || ((pixel_index >= 3769) && (pixel_index <= 3778)) || ((pixel_index >= 3793) && (pixel_index <= 3799)) || ((pixel_index >= 3864) && (pixel_index <= 3871)) || pixel_index == 3882 || ((pixel_index >= 3889) && (pixel_index <= 3897)) || ((pixel_index >= 3962) && (pixel_index <= 3964)) || pixel_index == 3978 || ((pixel_index >= 3985) && (pixel_index <= 3996)) || ((pixel_index >= 4059) && (pixel_index <= 4060)) || ((pixel_index >= 4074) && (pixel_index <= 4075)) || ((pixel_index >= 4081) && (pixel_index <= 4092)) || ((pixel_index >= 4155) && (pixel_index <= 4158)) || ((pixel_index >= 4170) && (pixel_index <= 4172)) || ((pixel_index >= 4177) && (pixel_index <= 4188)) || ((pixel_index >= 4251) && (pixel_index <= 4255)) || ((pixel_index >= 4266) && (pixel_index <= 4269)) || ((pixel_index >= 4274) && (pixel_index <= 4284)) || ((pixel_index >= 4347) && (pixel_index <= 4352)) || ((pixel_index >= 4362) && (pixel_index <= 4365)) || ((pixel_index >= 4370) && (pixel_index <= 4379)) || ((pixel_index >= 4444) && (pixel_index <= 4450)) || ((pixel_index >= 4459) && (pixel_index <= 4462)) || ((pixel_index >= 4467) && (pixel_index <= 4475)) || ((pixel_index >= 4480) && (pixel_index <= 4481)) || ((pixel_index >= 4541) && (pixel_index <= 4547)) || ((pixel_index >= 4555) && (pixel_index <= 4559)) || ((pixel_index >= 4575) && (pixel_index <= 4578)) || ((pixel_index >= 4637) && (pixel_index <= 4644)) || ((pixel_index >= 4651) && (pixel_index <= 4656)) || ((pixel_index >= 4670) && (pixel_index <= 4675)) || ((pixel_index >= 4677) && (pixel_index <= 4678)) || ((pixel_index >= 4734) && (pixel_index <= 4742)) || ((pixel_index >= 4747) && (pixel_index <= 4754)) || ((pixel_index >= 4766) && (pixel_index <= 4773)) || ((pixel_index >= 4831) && (pixel_index <= 4839)) || ((pixel_index >= 4844) && (pixel_index <= 4856)) || ((pixel_index >= 4861) && (pixel_index <= 4869)) || ((pixel_index >= 4928) && (pixel_index <= 4937)) || ((pixel_index >= 4940) && (pixel_index <= 4951)) || ((pixel_index >= 4956) && (pixel_index <= 4966)) || ((pixel_index >= 5026) && (pixel_index <= 5046)) || ((pixel_index >= 5051) && (pixel_index <= 5063)) || ((pixel_index >= 5122) && (pixel_index <= 5131)) || ((pixel_index >= 5133) && (pixel_index <= 5143)) || ((pixel_index >= 5145) && (pixel_index <= 5161)) || ((pixel_index >= 5218) && (pixel_index <= 5227)) || ((pixel_index >= 5229) && (pixel_index <= 5258)) || ((pixel_index >= 5314) && (pixel_index <= 5324)) || ((pixel_index >= 5326) && (pixel_index <= 5355)) || ((pixel_index >= 5410) && (pixel_index <= 5419)) || ((pixel_index >= 5422) && (pixel_index <= 5447)) || ((pixel_index >= 5450) && (pixel_index <= 5451)) || ((pixel_index >= 5505) && (pixel_index <= 5516)) || ((pixel_index >= 5519) && (pixel_index <= 5542)) || ((pixel_index >= 5546) && (pixel_index <= 5547)) || ((pixel_index >= 5602) && (pixel_index <= 5613)) || ((pixel_index >= 5615) && (pixel_index <= 5636)) || ((pixel_index >= 5640) && (pixel_index <= 5643)) || ((pixel_index >= 5699) && (pixel_index <= 5723)) || ((pixel_index >= 5727) && (pixel_index <= 5738)) || ((pixel_index >= 5794) && (pixel_index <= 5818)) || ((pixel_index >= 5825) && (pixel_index <= 5833)) || ((pixel_index >= 5891) && (pixel_index <= 5905)) || ((pixel_index >= 5909) && (pixel_index <= 5911)) || ((pixel_index >= 5925) && (pixel_index <= 5927)) || ((pixel_index >= 5987) && (pixel_index <= 6001)) || pixel_index == 6006 || (pixel_index >= 6085) && (pixel_index <= 6097)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 28) begin
            if (((pixel_index >= 2232) && (pixel_index <= 2235)) || ((pixel_index >= 2327) && (pixel_index <= 2333)) || ((pixel_index >= 2424) && (pixel_index <= 2430)) || ((pixel_index >= 2522) && (pixel_index <= 2527)) || ((pixel_index >= 2619) && (pixel_index <= 2624)) || ((pixel_index >= 2716) && (pixel_index <= 2720)) || ((pixel_index >= 2812) && (pixel_index <= 2817)) || ((pixel_index >= 2909) && (pixel_index <= 2913)) || pixel_index == 3009 || ((pixel_index >= 3412) && (pixel_index <= 3413)) || ((pixel_index >= 3508) && (pixel_index <= 3510)) || ((pixel_index >= 3575) && (pixel_index <= 3576)) || ((pixel_index >= 3604) && (pixel_index <= 3607)) || ((pixel_index >= 3671) && (pixel_index <= 3672)) || ((pixel_index >= 3700) && (pixel_index <= 3705)) || ((pixel_index >= 3766) && (pixel_index <= 3768)) || ((pixel_index >= 3796) && (pixel_index <= 3804)) || ((pixel_index >= 3862) && (pixel_index <= 3864)) || pixel_index == 3887 || ((pixel_index >= 3892) && (pixel_index <= 3902)) || ((pixel_index >= 3959) && (pixel_index <= 3961)) || pixel_index == 3983 || ((pixel_index >= 3989) && (pixel_index <= 3998)) || ((pixel_index >= 4055) && (pixel_index <= 4057)) || pixel_index == 4060 || ((pixel_index >= 4079) && (pixel_index <= 4080)) || ((pixel_index >= 4087) && (pixel_index <= 4094)) || ((pixel_index >= 4151) && (pixel_index <= 4154)) || ((pixel_index >= 4156) && (pixel_index <= 4157)) || ((pixel_index >= 4175) && (pixel_index <= 4176)) || ((pixel_index >= 4186) && (pixel_index <= 4189)) || ((pixel_index >= 4248) && (pixel_index <= 4251)) || ((pixel_index >= 4253) && (pixel_index <= 4254)) || ((pixel_index >= 4271) && (pixel_index <= 4273)) || ((pixel_index >= 4344) && (pixel_index <= 4352)) || ((pixel_index >= 4367) && (pixel_index <= 4369)) || ((pixel_index >= 4441) && (pixel_index <= 4449)) || ((pixel_index >= 4463) && (pixel_index <= 4466)) || ((pixel_index >= 4483) && (pixel_index <= 4484)) || pixel_index == 4490 || ((pixel_index >= 4538) && (pixel_index <= 4547)) || ((pixel_index >= 4559) && (pixel_index <= 4563)) || ((pixel_index >= 4578) && (pixel_index <= 4585)) || ((pixel_index >= 4635) && (pixel_index <= 4645)) || ((pixel_index >= 4655) && (pixel_index <= 4664)) || ((pixel_index >= 4673) && (pixel_index <= 4680)) || ((pixel_index >= 4732) && (pixel_index <= 4742)) || ((pixel_index >= 4751) && (pixel_index <= 4761)) || pixel_index == 4765 || ((pixel_index >= 4767) && (pixel_index <= 4775)) || ((pixel_index >= 4829) && (pixel_index <= 4841)) || ((pixel_index >= 4847) && (pixel_index <= 4856)) || ((pixel_index >= 4861) && (pixel_index <= 4871)) || ((pixel_index >= 4927) && (pixel_index <= 4938)) || ((pixel_index >= 4943) && (pixel_index <= 4951)) || ((pixel_index >= 4958) && (pixel_index <= 4967)) || ((pixel_index >= 5025) && (pixel_index <= 5034)) || ((pixel_index >= 5040) && (pixel_index <= 5047)) || ((pixel_index >= 5053) && (pixel_index <= 5064)) || ((pixel_index >= 5121) && (pixel_index <= 5130)) || ((pixel_index >= 5136) && (pixel_index <= 5144)) || ((pixel_index >= 5148) && (pixel_index <= 5162)) || ((pixel_index >= 5217) && (pixel_index <= 5226)) || ((pixel_index >= 5231) && (pixel_index <= 5240)) || ((pixel_index >= 5243) && (pixel_index <= 5259)) || ((pixel_index >= 5312) && (pixel_index <= 5323)) || ((pixel_index >= 5327) && (pixel_index <= 5356)) || ((pixel_index >= 5409) && (pixel_index <= 5420)) || ((pixel_index >= 5424) && (pixel_index <= 5453)) || ((pixel_index >= 5506) && (pixel_index <= 5517)) || ((pixel_index >= 5520) && (pixel_index <= 5549)) || ((pixel_index >= 5603) && (pixel_index <= 5616)) || ((pixel_index >= 5618) && (pixel_index <= 5630)) || ((pixel_index >= 5634) && (pixel_index <= 5645)) || ((pixel_index >= 5698) && (pixel_index <= 5712)) || ((pixel_index >= 5715) && (pixel_index <= 5727)) || ((pixel_index >= 5731) && (pixel_index <= 5733)) || ((pixel_index >= 5739) && (pixel_index <= 5741)) || ((pixel_index >= 5794) && (pixel_index <= 5808)) || ((pixel_index >= 5812) && (pixel_index <= 5822)) || ((pixel_index >= 5828) && (pixel_index <= 5831)) || ((pixel_index >= 5833) && (pixel_index <= 5836)) || ((pixel_index >= 5891) && (pixel_index <= 5905)) || ((pixel_index >= 5911) && (pixel_index <= 5917)) || ((pixel_index >= 5925) && (pixel_index <= 5931)) || ((pixel_index >= 5987) && (pixel_index <= 6001)) || pixel_index == 6010 || ((pixel_index >= 6024) && (pixel_index <= 6025)) || (pixel_index >= 6085) && (pixel_index <= 6095)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 29) begin
            if (((pixel_index >= 687) && (pixel_index <= 689)) || ((pixel_index >= 782) && (pixel_index <= 787)) || ((pixel_index >= 878) && (pixel_index <= 886)) || ((pixel_index >= 974) && (pixel_index <= 984)) || ((pixel_index >= 1070) && (pixel_index <= 1081)) || ((pixel_index >= 1167) && (pixel_index <= 1176)) || ((pixel_index >= 1263) && (pixel_index <= 1272)) || ((pixel_index >= 1360) && (pixel_index <= 1368)) || ((pixel_index >= 1457) && (pixel_index <= 1464)) || ((pixel_index >= 1554) && (pixel_index <= 1560)) || ((pixel_index >= 1651) && (pixel_index <= 1656)) || ((pixel_index >= 1748) && (pixel_index <= 1752)) || ((pixel_index >= 1845) && (pixel_index <= 1848)) || ((pixel_index >= 1942) && (pixel_index <= 1945)) || ((pixel_index >= 2039) && (pixel_index <= 2041)) || ((pixel_index >= 2136) && (pixel_index <= 2137)) || ((pixel_index >= 3318) && (pixel_index <= 3319)) || ((pixel_index >= 3414) && (pixel_index <= 3416)) || ((pixel_index >= 3510) && (pixel_index <= 3513)) || ((pixel_index >= 3570) && (pixel_index <= 3571)) || ((pixel_index >= 3607) && (pixel_index <= 3611)) || ((pixel_index >= 3666) && (pixel_index <= 3667)) || ((pixel_index >= 3704) && (pixel_index <= 3710)) || ((pixel_index >= 3762) && (pixel_index <= 3764)) || ((pixel_index >= 3802) && (pixel_index <= 3807)) || ((pixel_index >= 3858) && (pixel_index <= 3861)) || pixel_index == 3892 || ((pixel_index >= 3900) && (pixel_index <= 3903)) || ((pixel_index >= 3954) && (pixel_index <= 3957)) || pixel_index == 3962 || ((pixel_index >= 3988) && (pixel_index <= 3989)) || ((pixel_index >= 4051) && (pixel_index <= 4054)) || ((pixel_index >= 4058) && (pixel_index <= 4059)) || ((pixel_index >= 4084) && (pixel_index <= 4085)) || ((pixel_index >= 4147) && (pixel_index <= 4151)) || ((pixel_index >= 4155) && (pixel_index <= 4156)) || ((pixel_index >= 4180) && (pixel_index <= 4181)) || ((pixel_index >= 4244) && (pixel_index <= 4249)) || ((pixel_index >= 4252) && (pixel_index <= 4254)) || ((pixel_index >= 4276) && (pixel_index <= 4277)) || ((pixel_index >= 4295) && (pixel_index <= 4296)) || pixel_index == 4302 || ((pixel_index >= 4341) && (pixel_index <= 4351)) || ((pixel_index >= 4371) && (pixel_index <= 4374)) || ((pixel_index >= 4389) && (pixel_index <= 4394)) || ((pixel_index >= 4396) && (pixel_index <= 4398)) || ((pixel_index >= 4438) && (pixel_index <= 4449)) || ((pixel_index >= 4467) && (pixel_index <= 4470)) || ((pixel_index >= 4480) && (pixel_index <= 4493)) || ((pixel_index >= 4535) && (pixel_index <= 4548)) || ((pixel_index >= 4562) && (pixel_index <= 4568)) || ((pixel_index >= 4577) && (pixel_index <= 4586)) || ((pixel_index >= 4632) && (pixel_index <= 4646)) || ((pixel_index >= 4658) && (pixel_index <= 4666)) || ((pixel_index >= 4676) && (pixel_index <= 4678)) || ((pixel_index >= 4730) && (pixel_index <= 4744)) || ((pixel_index >= 4754) && (pixel_index <= 4761)) || ((pixel_index >= 4771) && (pixel_index <= 4774)) || ((pixel_index >= 4828) && (pixel_index <= 4841)) || ((pixel_index >= 4849) && (pixel_index <= 4856)) || ((pixel_index >= 4866) && (pixel_index <= 4871)) || ((pixel_index >= 4927) && (pixel_index <= 4937)) || ((pixel_index >= 4945) && (pixel_index <= 4952)) || ((pixel_index >= 4961) && (pixel_index <= 4968)) || ((pixel_index >= 5023) && (pixel_index <= 5033)) || ((pixel_index >= 5040) && (pixel_index <= 5049)) || ((pixel_index >= 5056) && (pixel_index <= 5065)) || ((pixel_index >= 5119) && (pixel_index <= 5129)) || ((pixel_index >= 5136) && (pixel_index <= 5145)) || ((pixel_index >= 5150) && (pixel_index <= 5161)) || ((pixel_index >= 5216) && (pixel_index <= 5227)) || ((pixel_index >= 5233) && (pixel_index <= 5242)) || ((pixel_index >= 5245) && (pixel_index <= 5258)) || ((pixel_index >= 5313) && (pixel_index <= 5321)) || ((pixel_index >= 5330) && (pixel_index <= 5356)) || ((pixel_index >= 5409) && (pixel_index <= 5423)) || ((pixel_index >= 5427) && (pixel_index <= 5453)) || ((pixel_index >= 5506) && (pixel_index <= 5519)) || ((pixel_index >= 5523) && (pixel_index <= 5532)) || ((pixel_index >= 5534) && (pixel_index <= 5536)) || ((pixel_index >= 5540) && (pixel_index <= 5550)) || ((pixel_index >= 5602) && (pixel_index <= 5615)) || ((pixel_index >= 5620) && (pixel_index <= 5629)) || ((pixel_index >= 5637) && (pixel_index <= 5638)) || ((pixel_index >= 5641) && (pixel_index <= 5646)) || ((pixel_index >= 5698) && (pixel_index <= 5712)) || ((pixel_index >= 5716) && (pixel_index <= 5726)) || ((pixel_index >= 5733) && (pixel_index <= 5734)) || ((pixel_index >= 5738) && (pixel_index <= 5742)) || ((pixel_index >= 5794) && (pixel_index <= 5808)) || ((pixel_index >= 5814) && (pixel_index <= 5823)) || ((pixel_index >= 5830) && (pixel_index <= 5831)) || ((pixel_index >= 5836) && (pixel_index <= 5837)) || ((pixel_index >= 5890) && (pixel_index <= 5904)) || ((pixel_index >= 5911) && (pixel_index <= 5920)) || ((pixel_index >= 5926) && (pixel_index <= 5928)) || ((pixel_index >= 5930) && (pixel_index <= 5933)) || ((pixel_index >= 5987) && (pixel_index <= 5998)) || ((pixel_index >= 6009) && (pixel_index <= 6016)) || ((pixel_index >= 6024) && (pixel_index <= 6028)) || ((pixel_index >= 6085) && (pixel_index <= 6091)) || ((pixel_index >= 6107) && (pixel_index <= 6110)) || (pixel_index >= 6121) && (pixel_index <= 6123)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 30) begin
            if (pixel_index == 309 || ((pixel_index >= 404) && (pixel_index <= 405)) || pixel_index == 500 || ((pixel_index >= 595) && (pixel_index <= 596)) || ((pixel_index >= 690) && (pixel_index <= 692)) || ((pixel_index >= 785) && (pixel_index <= 787)) || ((pixel_index >= 879) && (pixel_index <= 883)) || ((pixel_index >= 970) && (pixel_index <= 978)) || ((pixel_index >= 1065) && (pixel_index <= 1074)) || ((pixel_index >= 1160) && (pixel_index <= 1169)) || ((pixel_index >= 1257) && (pixel_index <= 1264)) || ((pixel_index >= 1354) && (pixel_index <= 1358)) || ((pixel_index >= 3320) && (pixel_index <= 3321)) || ((pixel_index >= 3417) && (pixel_index <= 3418)) || ((pixel_index >= 3513) && (pixel_index <= 3517)) || ((pixel_index >= 3610) && (pixel_index <= 3614)) || ((pixel_index >= 3707) && (pixel_index <= 3711)) || pixel_index == 3761 || ((pixel_index >= 3805) && (pixel_index <= 3809)) || ((pixel_index >= 3857) && (pixel_index <= 3858)) || ((pixel_index >= 3903) && (pixel_index <= 3906)) || ((pixel_index >= 3952) && (pixel_index <= 3955)) || ((pixel_index >= 4049) && (pixel_index <= 4051)) || pixel_index == 4058 || pixel_index == 4090 || ((pixel_index >= 4145) && (pixel_index <= 4148)) || ((pixel_index >= 4154) && (pixel_index <= 4155)) || pixel_index == 4186 || ((pixel_index >= 4241) && (pixel_index <= 4246)) || ((pixel_index >= 4251) && (pixel_index <= 4252)) || ((pixel_index >= 4281) && (pixel_index <= 4282)) || ((pixel_index >= 4299) && (pixel_index <= 4300)) || ((pixel_index >= 4338) && (pixel_index <= 4345)) || ((pixel_index >= 4347) && (pixel_index <= 4350)) || ((pixel_index >= 4377) && (pixel_index <= 4378)) || ((pixel_index >= 4388) && (pixel_index <= 4390)) || ((pixel_index >= 4393) && (pixel_index <= 4398)) || ((pixel_index >= 4402) && (pixel_index <= 4403)) || ((pixel_index >= 4435) && (pixel_index <= 4448)) || pixel_index == 4469 || ((pixel_index >= 4473) && (pixel_index <= 4475)) || ((pixel_index >= 4485) && (pixel_index <= 4499)) || ((pixel_index >= 4532) && (pixel_index <= 4546)) || ((pixel_index >= 4564) && (pixel_index <= 4571)) || ((pixel_index >= 4583) && (pixel_index <= 4594)) || ((pixel_index >= 4629) && (pixel_index <= 4645)) || ((pixel_index >= 4660) && (pixel_index <= 4668)) || ((pixel_index >= 4682) && (pixel_index <= 4687)) || ((pixel_index >= 4726) && (pixel_index <= 4744)) || ((pixel_index >= 4755) && (pixel_index <= 4765)) || ((pixel_index >= 4823) && (pixel_index <= 4841)) || ((pixel_index >= 4851) && (pixel_index <= 4860)) || ((pixel_index >= 4870) && (pixel_index <= 4872)) || ((pixel_index >= 4921) && (pixel_index <= 4938)) || ((pixel_index >= 4946) && (pixel_index <= 4956)) || ((pixel_index >= 4965) && (pixel_index <= 4969)) || ((pixel_index >= 5020) && (pixel_index <= 5034)) || ((pixel_index >= 5042) && (pixel_index <= 5052)) || ((pixel_index >= 5060) && (pixel_index <= 5065)) || ((pixel_index >= 5120) && (pixel_index <= 5130)) || ((pixel_index >= 5138) && (pixel_index <= 5148)) || ((pixel_index >= 5155) && (pixel_index <= 5162)) || ((pixel_index >= 5216) && (pixel_index <= 5228)) || ((pixel_index >= 5235) && (pixel_index <= 5245)) || ((pixel_index >= 5249) && (pixel_index <= 5258)) || ((pixel_index >= 5313) && (pixel_index <= 5322)) || ((pixel_index >= 5332) && (pixel_index <= 5341)) || ((pixel_index >= 5345) && (pixel_index <= 5355)) || ((pixel_index >= 5409) && (pixel_index <= 5416)) || ((pixel_index >= 5430) && (pixel_index <= 5437)) || ((pixel_index >= 5442) && (pixel_index <= 5452)) || ((pixel_index >= 5505) && (pixel_index <= 5520)) || ((pixel_index >= 5526) && (pixel_index <= 5534)) || ((pixel_index >= 5539) && (pixel_index <= 5551)) || ((pixel_index >= 5602) && (pixel_index <= 5616)) || ((pixel_index >= 5622) && (pixel_index <= 5630)) || ((pixel_index >= 5639) && (pixel_index <= 5648)) || ((pixel_index >= 5699) && (pixel_index <= 5713)) || ((pixel_index >= 5718) && (pixel_index <= 5727)) || ((pixel_index >= 5736) && (pixel_index <= 5744)) || ((pixel_index >= 5795) && (pixel_index <= 5809)) || ((pixel_index >= 5815) && (pixel_index <= 5823)) || ((pixel_index >= 5832) && (pixel_index <= 5833)) || ((pixel_index >= 5836) && (pixel_index <= 5841)) || ((pixel_index >= 5891) && (pixel_index <= 5906)) || ((pixel_index >= 5911) && (pixel_index <= 5920)) || ((pixel_index >= 5928) && (pixel_index <= 5929)) || ((pixel_index >= 5932) && (pixel_index <= 5936)) || ((pixel_index >= 5987) && (pixel_index <= 6001)) || ((pixel_index >= 6009) && (pixel_index <= 6016)) || ((pixel_index >= 6024) && (pixel_index <= 6026)) || ((pixel_index >= 6029) && (pixel_index <= 6032)) || ((pixel_index >= 6084) && (pixel_index <= 6096)) || ((pixel_index >= 6106) && (pixel_index <= 6113)) || ((pixel_index >= 6121) && (pixel_index <= 6122)) || (pixel_index >= 6125) && (pixel_index <= 6127)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 31) begin
            oled_data = 0;
            done = 1;
        end
    end
    
endmodule

module draw_anim(input frame_rate, input start, input [12:0] pixel_index, output reg done, output reg [15:0] oled_data);
    reg [15:0] frame_count = 0;
    
    always @ (posedge frame_rate) begin
        if (start) frame_count <= (frame_count == 31) ? 31 : frame_count + 1;
        else frame_count <= 0;
    end
   
    // animation for player draw (AI mode only)
    // Reimu and Marisa after yin yang
    always @ (*) begin
        if (frame_count <= 30) done = 0;
        if (frame_count == 0) oled_data = 0;
        else if (frame_count == 1) begin
            if (((pixel_index >= 5) && (pixel_index <= 47)) || ((pixel_index >= 79) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 144)) || ((pixel_index >= 176) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 240)) || ((pixel_index >= 273) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 337)) || ((pixel_index >= 370) && (pixel_index <= 377)) || ((pixel_index >= 389) && (pixel_index <= 394)) || ((pixel_index >= 396) && (pixel_index <= 434)) || ((pixel_index >= 467) && (pixel_index <= 473)) || ((pixel_index >= 485) && (pixel_index <= 489)) || ((pixel_index >= 491) && (pixel_index <= 530)) || ((pixel_index >= 564) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 584)) || ((pixel_index >= 586) && (pixel_index <= 627)) || ((pixel_index >= 660) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 679)) || ((pixel_index >= 682) && (pixel_index <= 723)) || ((pixel_index >= 757) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 774)) || ((pixel_index >= 777) && (pixel_index <= 820)) || ((pixel_index >= 853) && (pixel_index <= 857)) || pixel_index == 869 || ((pixel_index >= 873) && (pixel_index <= 916)) || ((pixel_index >= 950) && (pixel_index <= 953)) || ((pixel_index >= 968) && (pixel_index <= 1012)) || ((pixel_index >= 1047) && (pixel_index <= 1049)) || ((pixel_index >= 1064) && (pixel_index <= 1085)) || ((pixel_index >= 1091) && (pixel_index <= 1108)) || ((pixel_index >= 1143) && (pixel_index <= 1145)) || ((pixel_index >= 1159) && (pixel_index <= 1180)) || ((pixel_index >= 1189) && (pixel_index <= 1205)) || ((pixel_index >= 1240) && (pixel_index <= 1241)) || ((pixel_index >= 1254) && (pixel_index <= 1275)) || ((pixel_index >= 1286) && (pixel_index <= 1301)) || ((pixel_index >= 1336) && (pixel_index <= 1337)) || ((pixel_index >= 1350) && (pixel_index <= 1370)) || ((pixel_index >= 1382) && (pixel_index <= 1397)) || pixel_index == 1433 || ((pixel_index >= 1446) && (pixel_index <= 1466)) || ((pixel_index >= 1478) && (pixel_index <= 1493)) || pixel_index == 1529 || ((pixel_index >= 1541) && (pixel_index <= 1562)) || ((pixel_index >= 1574) && (pixel_index <= 1589)) || pixel_index == 1625 || ((pixel_index >= 1637) && (pixel_index <= 1658)) || ((pixel_index >= 1670) && (pixel_index <= 1685)) || ((pixel_index >= 1733) && (pixel_index <= 1754)) || ((pixel_index >= 1766) && (pixel_index <= 1781)) || ((pixel_index >= 1829) && (pixel_index <= 1850)) || ((pixel_index >= 1862) && (pixel_index <= 1877)) || ((pixel_index >= 1925) && (pixel_index <= 1947)) || ((pixel_index >= 1957) && (pixel_index <= 1972)) || ((pixel_index >= 2021) && (pixel_index <= 2044)) || ((pixel_index >= 2052) && (pixel_index <= 2068)) || ((pixel_index >= 2117) && (pixel_index <= 2142)) || ((pixel_index >= 2146) && (pixel_index <= 2164)) || ((pixel_index >= 2213) && (pixel_index <= 2260)) || ((pixel_index >= 2309) && (pixel_index <= 2355)) || ((pixel_index >= 2405) && (pixel_index <= 2451)) || ((pixel_index >= 2501) && (pixel_index <= 2546)) || ((pixel_index >= 2597) && (pixel_index <= 2642)) || ((pixel_index >= 2693) && (pixel_index <= 2737)) || ((pixel_index >= 2789) && (pixel_index <= 2833)) || ((pixel_index >= 2885) && (pixel_index <= 2928)) || ((pixel_index >= 2981) && (pixel_index <= 3023)) || ((pixel_index >= 3077) && (pixel_index <= 3118)) || ((pixel_index >= 3173) && (pixel_index <= 3213)) || ((pixel_index >= 3269) && (pixel_index <= 3308)) || ((pixel_index >= 3365) && (pixel_index <= 3403)) || ((pixel_index >= 3461) && (pixel_index <= 3499)) || ((pixel_index >= 3557) && (pixel_index <= 3594)) || ((pixel_index >= 3653) && (pixel_index <= 3690)) || ((pixel_index >= 3749) && (pixel_index <= 3785)) || ((pixel_index >= 3845) && (pixel_index <= 3881)) || ((pixel_index >= 3941) && (pixel_index <= 3977)) || ((pixel_index >= 4037) && (pixel_index <= 4072)) || ((pixel_index >= 4092) && (pixel_index <= 4096)) || ((pixel_index >= 4133) && (pixel_index <= 4168)) || ((pixel_index >= 4187) && (pixel_index <= 4194)) || ((pixel_index >= 4229) && (pixel_index <= 4264)) || ((pixel_index >= 4282) && (pixel_index <= 4290)) || ((pixel_index >= 4325) && (pixel_index <= 4360)) || ((pixel_index >= 4377) && (pixel_index <= 4387)) || ((pixel_index >= 4421) && (pixel_index <= 4456)) || ((pixel_index >= 4473) && (pixel_index <= 4483)) || ((pixel_index >= 4517) && (pixel_index <= 4552)) || ((pixel_index >= 4569) && (pixel_index <= 4579)) || pixel_index == 4601 || ((pixel_index >= 4614) && (pixel_index <= 4648)) || ((pixel_index >= 4665) && (pixel_index <= 4675)) || pixel_index == 4697 || ((pixel_index >= 4710) && (pixel_index <= 4744)) || ((pixel_index >= 4761) && (pixel_index <= 4770)) || pixel_index == 4793 || ((pixel_index >= 4807) && (pixel_index <= 4840)) || ((pixel_index >= 4858) && (pixel_index <= 4866)) || ((pixel_index >= 4888) && (pixel_index <= 4889)) || ((pixel_index >= 4903) && (pixel_index <= 4936)) || ((pixel_index >= 4955) && (pixel_index <= 4961)) || ((pixel_index >= 4984) && (pixel_index <= 4985)) || ((pixel_index >= 4999) && (pixel_index <= 5032)) || ((pixel_index >= 5053) && (pixel_index <= 5055)) || ((pixel_index >= 5079) && (pixel_index <= 5081)) || ((pixel_index >= 5096) && (pixel_index <= 5128)) || ((pixel_index >= 5175) && (pixel_index <= 5177)) || ((pixel_index >= 5193) && (pixel_index <= 5225)) || ((pixel_index >= 5270) && (pixel_index <= 5272)) || ((pixel_index >= 5289) && (pixel_index <= 5321)) || ((pixel_index >= 5365) && (pixel_index <= 5367)) || ((pixel_index >= 5386) && (pixel_index <= 5417)) || ((pixel_index >= 5461) && (pixel_index <= 5462)) || ((pixel_index >= 5482) && (pixel_index <= 5514)) || ((pixel_index >= 5556) && (pixel_index <= 5557)) || ((pixel_index >= 5579) && (pixel_index <= 5610)) || pixel_index == 5652 || ((pixel_index >= 5676) && (pixel_index <= 5707)) || pixel_index == 5747 || ((pixel_index >= 5773) && (pixel_index <= 5804)) || pixel_index == 5842 || ((pixel_index >= 5870) && (pixel_index <= 5900)) || ((pixel_index >= 5967) && (pixel_index <= 5997)) || (pixel_index >= 6063) && (pixel_index <= 6094)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 2) begin
            if (((pixel_index >= 14) && (pixel_index <= 79)) || ((pixel_index >= 81) && (pixel_index <= 89)) || ((pixel_index >= 109) && (pixel_index <= 176)) || ((pixel_index >= 178) && (pixel_index <= 185)) || ((pixel_index >= 204) && (pixel_index <= 272)) || ((pixel_index >= 275) && (pixel_index <= 281)) || ((pixel_index >= 299) && (pixel_index <= 369)) || ((pixel_index >= 372) && (pixel_index <= 377)) || ((pixel_index >= 395) && (pixel_index <= 465)) || ((pixel_index >= 468) && (pixel_index <= 473)) || ((pixel_index >= 490) && (pixel_index <= 562)) || ((pixel_index >= 565) && (pixel_index <= 569)) || ((pixel_index >= 585) && (pixel_index <= 658)) || ((pixel_index >= 662) && (pixel_index <= 665)) || ((pixel_index >= 680) && (pixel_index <= 754)) || ((pixel_index >= 758) && (pixel_index <= 761)) || ((pixel_index >= 776) && (pixel_index <= 851)) || ((pixel_index >= 855) && (pixel_index <= 857)) || ((pixel_index >= 871) && (pixel_index <= 921)) || ((pixel_index >= 928) && (pixel_index <= 947)) || ((pixel_index >= 952) && (pixel_index <= 953)) || ((pixel_index >= 967) && (pixel_index <= 1015)) || ((pixel_index >= 1025) && (pixel_index <= 1043)) || ((pixel_index >= 1048) && (pixel_index <= 1049)) || ((pixel_index >= 1062) && (pixel_index <= 1111)) || ((pixel_index >= 1122) && (pixel_index <= 1139)) || pixel_index == 1145 || ((pixel_index >= 1158) && (pixel_index <= 1206)) || ((pixel_index >= 1218) && (pixel_index <= 1235)) || pixel_index == 1241 || ((pixel_index >= 1253) && (pixel_index <= 1302)) || ((pixel_index >= 1314) && (pixel_index <= 1331)) || ((pixel_index >= 1349) && (pixel_index <= 1398)) || ((pixel_index >= 1410) && (pixel_index <= 1427)) || ((pixel_index >= 1445) && (pixel_index <= 1494)) || ((pixel_index >= 1506) && (pixel_index <= 1523)) || ((pixel_index >= 1541) && (pixel_index <= 1590)) || ((pixel_index >= 1602) && (pixel_index <= 1619)) || ((pixel_index >= 1637) && (pixel_index <= 1686)) || ((pixel_index >= 1698) && (pixel_index <= 1715)) || ((pixel_index >= 1733) && (pixel_index <= 1783)) || ((pixel_index >= 1793) && (pixel_index <= 1811)) || ((pixel_index >= 1829) && (pixel_index <= 1880)) || ((pixel_index >= 1888) && (pixel_index <= 1906)) || ((pixel_index >= 1925) && (pixel_index <= 1978)) || ((pixel_index >= 1982) && (pixel_index <= 2002)) || ((pixel_index >= 2021) && (pixel_index <= 2098)) || ((pixel_index >= 2117) && (pixel_index <= 2193)) || ((pixel_index >= 2213) && (pixel_index <= 2289)) || ((pixel_index >= 2309) && (pixel_index <= 2384)) || ((pixel_index >= 2405) && (pixel_index <= 2480)) || ((pixel_index >= 2501) && (pixel_index <= 2575)) || ((pixel_index >= 2597) && (pixel_index <= 2622)) || ((pixel_index >= 2629) && (pixel_index <= 2670)) || ((pixel_index >= 2693) && (pixel_index <= 2713)) || ((pixel_index >= 2729) && (pixel_index <= 2766)) || ((pixel_index >= 2789) && (pixel_index <= 2807)) || ((pixel_index >= 2828) && (pixel_index <= 2861)) || ((pixel_index >= 2885) && (pixel_index <= 2901)) || ((pixel_index >= 2926) && (pixel_index <= 2956)) || ((pixel_index >= 2981) && (pixel_index <= 2996)) || ((pixel_index >= 3023) && (pixel_index <= 3050)) || ((pixel_index >= 3077) && (pixel_index <= 3090)) || ((pixel_index >= 3120) && (pixel_index <= 3145)) || ((pixel_index >= 3173) && (pixel_index <= 3185)) || ((pixel_index >= 3218) && (pixel_index <= 3240)) || ((pixel_index >= 3269) && (pixel_index <= 3280)) || ((pixel_index >= 3316) && (pixel_index <= 3334)) || ((pixel_index >= 3365) && (pixel_index <= 3375)) || ((pixel_index >= 3415) && (pixel_index <= 3427)) || ((pixel_index >= 3461) && (pixel_index <= 3470)) || ((pixel_index >= 3516) && (pixel_index <= 3518)) || ((pixel_index >= 3557) && (pixel_index <= 3565)) || ((pixel_index >= 3653) && (pixel_index <= 3661)) || ((pixel_index >= 3749) && (pixel_index <= 3756)) || ((pixel_index >= 3845) && (pixel_index <= 3852)) || ((pixel_index >= 3941) && (pixel_index <= 3947)) || ((pixel_index >= 4037) && (pixel_index <= 4043)) || ((pixel_index >= 4133) && (pixel_index <= 4139)) || ((pixel_index >= 4229) && (pixel_index <= 4235)) || ((pixel_index >= 4255) && (pixel_index <= 4260)) || ((pixel_index >= 4325) && (pixel_index <= 4330)) || ((pixel_index >= 4350) && (pixel_index <= 4357)) || ((pixel_index >= 4421) && (pixel_index <= 4426)) || ((pixel_index >= 4445) && (pixel_index <= 4454)) || ((pixel_index >= 4517) && (pixel_index <= 4522)) || ((pixel_index >= 4541) && (pixel_index <= 4551)) || ((pixel_index >= 4613) && (pixel_index <= 4618)) || ((pixel_index >= 4637) && (pixel_index <= 4647)) || ((pixel_index >= 4709) && (pixel_index <= 4714)) || ((pixel_index >= 4733) && (pixel_index <= 4743)) || ((pixel_index >= 4805) && (pixel_index <= 4810)) || ((pixel_index >= 4829) && (pixel_index <= 4839)) || ((pixel_index >= 4902) && (pixel_index <= 4906)) || ((pixel_index >= 4925) && (pixel_index <= 4935)) || pixel_index == 4985 || ((pixel_index >= 4998) && (pixel_index <= 5002)) || ((pixel_index >= 5022) && (pixel_index <= 5030)) || ((pixel_index >= 5080) && (pixel_index <= 5081)) || ((pixel_index >= 5095) && (pixel_index <= 5098)) || ((pixel_index >= 5119) && (pixel_index <= 5125)) || ((pixel_index >= 5176) && (pixel_index <= 5177)) || ((pixel_index >= 5191) && (pixel_index <= 5194)) || ((pixel_index >= 5216) && (pixel_index <= 5220)) || ((pixel_index >= 5271) && (pixel_index <= 5273)) || ((pixel_index >= 5288) && (pixel_index <= 5290)) || ((pixel_index >= 5367) && (pixel_index <= 5369)) || ((pixel_index >= 5385) && (pixel_index <= 5387)) || ((pixel_index >= 5462) && (pixel_index <= 5465)) || ((pixel_index >= 5481) && (pixel_index <= 5483)) || ((pixel_index >= 5558) && (pixel_index <= 5561)) || ((pixel_index >= 5578) && (pixel_index <= 5579)) || ((pixel_index >= 5653) && (pixel_index <= 5657)) || ((pixel_index >= 5675) && (pixel_index <= 5676)) || ((pixel_index >= 5748) && (pixel_index <= 5753)) || ((pixel_index >= 5771) && (pixel_index <= 5772)) || ((pixel_index >= 5844) && (pixel_index <= 5849)) || ((pixel_index >= 5868) && (pixel_index <= 5869)) || ((pixel_index >= 5939) && (pixel_index <= 5945)) || ((pixel_index >= 6034) && (pixel_index <= 6041)) || (pixel_index >= 6129) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 3) begin
            if (pixel_index == 13 || ((pixel_index >= 40) && (pixel_index <= 82)) || pixel_index == 108 || ((pixel_index >= 137) && (pixel_index <= 179)) || ((pixel_index >= 235) && (pixel_index <= 276)) || ((pixel_index >= 332) && (pixel_index <= 372)) || ((pixel_index >= 429) && (pixel_index <= 469)) || ((pixel_index >= 526) && (pixel_index <= 566)) || ((pixel_index >= 622) && (pixel_index <= 662)) || ((pixel_index >= 719) && (pixel_index <= 759)) || ((pixel_index >= 816) && (pixel_index <= 856)) || ((pixel_index >= 912) && (pixel_index <= 952)) || ((pixel_index >= 1009) && (pixel_index <= 1049)) || ((pixel_index >= 1105) && (pixel_index <= 1145)) || ((pixel_index >= 1201) && (pixel_index <= 1241)) || ((pixel_index >= 1298) && (pixel_index <= 1337)) || ((pixel_index >= 1394) && (pixel_index <= 1433)) || ((pixel_index >= 1466) && (pixel_index <= 1471)) || ((pixel_index >= 1490) && (pixel_index <= 1529)) || ((pixel_index >= 1561) && (pixel_index <= 1568)) || ((pixel_index >= 1586) && (pixel_index <= 1625)) || ((pixel_index >= 1656) && (pixel_index <= 1664)) || ((pixel_index >= 1683) && (pixel_index <= 1721)) || ((pixel_index >= 1751) && (pixel_index <= 1761)) || ((pixel_index >= 1779) && (pixel_index <= 1817)) || ((pixel_index >= 1847) && (pixel_index <= 1857)) || ((pixel_index >= 1875) && (pixel_index <= 1913)) || ((pixel_index >= 1943) && (pixel_index <= 1953)) || ((pixel_index >= 1971) && (pixel_index <= 2009)) || ((pixel_index >= 2039) && (pixel_index <= 2049)) || ((pixel_index >= 2067) && (pixel_index <= 2105)) || ((pixel_index >= 2135) && (pixel_index <= 2145)) || ((pixel_index >= 2163) && (pixel_index <= 2201)) || ((pixel_index >= 2231) && (pixel_index <= 2240)) || ((pixel_index >= 2259) && (pixel_index <= 2297)) || ((pixel_index >= 2328) && (pixel_index <= 2335)) || ((pixel_index >= 2354) && (pixel_index <= 2393)) || ((pixel_index >= 2425) && (pixel_index <= 2430)) || ((pixel_index >= 2450) && (pixel_index <= 2489)) || ((pixel_index >= 2546) && (pixel_index <= 2585)) || ((pixel_index >= 2642) && (pixel_index <= 2681)) || ((pixel_index >= 2737) && (pixel_index <= 2777)) || ((pixel_index >= 2833) && (pixel_index <= 2873)) || ((pixel_index >= 2928) && (pixel_index <= 2969)) || ((pixel_index >= 3024) && (pixel_index <= 3065)) || ((pixel_index >= 3119) && (pixel_index <= 3161)) || ((pixel_index >= 3215) && (pixel_index <= 3257)) || ((pixel_index >= 3310) && (pixel_index <= 3353)) || ((pixel_index >= 3406) && (pixel_index <= 3449)) || ((pixel_index >= 3502) && (pixel_index <= 3545)) || ((pixel_index >= 3597) && (pixel_index <= 3616)) || ((pixel_index >= 3621) && (pixel_index <= 3641)) || ((pixel_index >= 3693) && (pixel_index <= 3710)) || ((pixel_index >= 3718) && (pixel_index <= 3737)) || ((pixel_index >= 3789) && (pixel_index <= 3805)) || ((pixel_index >= 3816) && (pixel_index <= 3833)) || ((pixel_index >= 3885) && (pixel_index <= 3900)) || ((pixel_index >= 3912) && (pixel_index <= 3929)) || ((pixel_index >= 3981) && (pixel_index <= 3996)) || ((pixel_index >= 4008) && (pixel_index <= 4025)) || ((pixel_index >= 4077) && (pixel_index <= 4092)) || ((pixel_index >= 4105) && (pixel_index <= 4121)) || ((pixel_index >= 4173) && (pixel_index <= 4187)) || ((pixel_index >= 4201) && (pixel_index <= 4217)) || ((pixel_index >= 4269) && (pixel_index <= 4284)) || ((pixel_index >= 4297) && (pixel_index <= 4313)) || ((pixel_index >= 4365) && (pixel_index <= 4380)) || ((pixel_index >= 4392) && (pixel_index <= 4409)) || ((pixel_index >= 4461) && (pixel_index <= 4476)) || ((pixel_index >= 4488) && (pixel_index <= 4505)) || ((pixel_index >= 4557) && (pixel_index <= 4573)) || ((pixel_index >= 4583) && (pixel_index <= 4601)) || ((pixel_index >= 4653) && (pixel_index <= 4670)) || ((pixel_index >= 4678) && (pixel_index <= 4697)) || ((pixel_index >= 4749) && (pixel_index <= 4768)) || ((pixel_index >= 4772) && (pixel_index <= 4793)) || ((pixel_index >= 4845) && (pixel_index <= 4889)) || ((pixel_index >= 4942) && (pixel_index <= 4985)) || ((pixel_index >= 5038) && (pixel_index <= 5081)) || pixel_index == 5093 || ((pixel_index >= 5134) && (pixel_index <= 5177)) || pixel_index == 5189 || ((pixel_index >= 5231) && (pixel_index <= 5273)) || ((pixel_index >= 5285) && (pixel_index <= 5286)) || ((pixel_index >= 5328) && (pixel_index <= 5369)) || ((pixel_index >= 5381) && (pixel_index <= 5382)) || ((pixel_index >= 5424) && (pixel_index <= 5465)) || ((pixel_index >= 5477) && (pixel_index <= 5479)) || ((pixel_index >= 5521) && (pixel_index <= 5561)) || ((pixel_index >= 5573) && (pixel_index <= 5576)) || ((pixel_index >= 5618) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5672)) || ((pixel_index >= 5714) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5769)) || ((pixel_index >= 5811) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5866)) || ((pixel_index >= 5908) && (pixel_index <= 5938)) || ((pixel_index >= 5940) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 5963)) || ((pixel_index >= 6006) && (pixel_index <= 6033)) || ((pixel_index >= 6035) && (pixel_index <= 6041)) || ((pixel_index >= 6053) && (pixel_index <= 6060)) || ((pixel_index >= 6103) && (pixel_index <= 6128)) || (pixel_index >= 6131) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 4) begin
            if (((pixel_index >= 5) && (pixel_index <= 10)) || ((pixel_index >= 80) && (pixel_index <= 83)) || ((pixel_index >= 101) && (pixel_index <= 105)) || ((pixel_index >= 176) && (pixel_index <= 180)) || ((pixel_index >= 197) && (pixel_index <= 200)) || ((pixel_index >= 273) && (pixel_index <= 277)) || ((pixel_index >= 293) && (pixel_index <= 296)) || ((pixel_index >= 369) && (pixel_index <= 374)) || ((pixel_index >= 389) && (pixel_index <= 391)) || ((pixel_index >= 465) && (pixel_index <= 470)) || ((pixel_index >= 485) && (pixel_index <= 486)) || ((pixel_index >= 561) && (pixel_index <= 567)) || ((pixel_index >= 581) && (pixel_index <= 582)) || ((pixel_index >= 630) && (pixel_index <= 635)) || ((pixel_index >= 657) && (pixel_index <= 664)) || pixel_index == 677 || ((pixel_index >= 725) && (pixel_index <= 733)) || ((pixel_index >= 754) && (pixel_index <= 760)) || ((pixel_index >= 820) && (pixel_index <= 829)) || ((pixel_index >= 850) && (pixel_index <= 857)) || ((pixel_index >= 916) && (pixel_index <= 926)) || ((pixel_index >= 946) && (pixel_index <= 953)) || ((pixel_index >= 1011) && (pixel_index <= 1022)) || ((pixel_index >= 1042) && (pixel_index <= 1049)) || ((pixel_index >= 1107) && (pixel_index <= 1118)) || ((pixel_index >= 1138) && (pixel_index <= 1145)) || ((pixel_index >= 1203) && (pixel_index <= 1214)) || ((pixel_index >= 1234) && (pixel_index <= 1241)) || ((pixel_index >= 1300) && (pixel_index <= 1310)) || ((pixel_index >= 1329) && (pixel_index <= 1337)) || ((pixel_index >= 1396) && (pixel_index <= 1405)) || ((pixel_index >= 1425) && (pixel_index <= 1433)) || ((pixel_index >= 1493) && (pixel_index <= 1501)) || ((pixel_index >= 1521) && (pixel_index <= 1529)) || ((pixel_index >= 1591) && (pixel_index <= 1595)) || ((pixel_index >= 1617) && (pixel_index <= 1625)) || ((pixel_index >= 1713) && (pixel_index <= 1721)) || ((pixel_index >= 1808) && (pixel_index <= 1817)) || ((pixel_index >= 1904) && (pixel_index <= 1913)) || ((pixel_index >= 1999) && (pixel_index <= 2009)) || ((pixel_index >= 2095) && (pixel_index <= 2105)) || ((pixel_index >= 2190) && (pixel_index <= 2201)) || ((pixel_index >= 2286) && (pixel_index <= 2297)) || ((pixel_index >= 2381) && (pixel_index <= 2393)) || ((pixel_index >= 2476) && (pixel_index <= 2489)) || ((pixel_index >= 2571) && (pixel_index <= 2585)) || ((pixel_index >= 2666) && (pixel_index <= 2681)) || ((pixel_index >= 2761) && (pixel_index <= 2777)) || ((pixel_index >= 2856) && (pixel_index <= 2873)) || ((pixel_index >= 2912) && (pixel_index <= 2921)) || ((pixel_index >= 2950) && (pixel_index <= 2969)) || ((pixel_index >= 3005) && (pixel_index <= 3021)) || ((pixel_index >= 3045) && (pixel_index <= 3065)) || ((pixel_index >= 3099) && (pixel_index <= 3119)) || ((pixel_index >= 3138) && (pixel_index <= 3161)) || ((pixel_index >= 3193) && (pixel_index <= 3218)) || ((pixel_index >= 3231) && (pixel_index <= 3257)) || ((pixel_index >= 3287) && (pixel_index <= 3353)) || ((pixel_index >= 3382) && (pixel_index <= 3449)) || ((pixel_index >= 3477) && (pixel_index <= 3545)) || ((pixel_index >= 3572) && (pixel_index <= 3641)) || ((pixel_index >= 3667) && (pixel_index <= 3737)) || ((pixel_index >= 3762) && (pixel_index <= 3833)) || ((pixel_index >= 3858) && (pixel_index <= 3929)) || ((pixel_index >= 3953) && (pixel_index <= 4025)) || ((pixel_index >= 4048) && (pixel_index <= 4121)) || ((pixel_index >= 4144) && (pixel_index <= 4217)) || ((pixel_index >= 4239) && (pixel_index <= 4313)) || ((pixel_index >= 4335) && (pixel_index <= 4409)) || ((pixel_index >= 4431) && (pixel_index <= 4451)) || ((pixel_index >= 4456) && (pixel_index <= 4505)) || ((pixel_index >= 4526) && (pixel_index <= 4545)) || ((pixel_index >= 4554) && (pixel_index <= 4601)) || ((pixel_index >= 4622) && (pixel_index <= 4640)) || ((pixel_index >= 4651) && (pixel_index <= 4697)) || ((pixel_index >= 4718) && (pixel_index <= 4735)) || ((pixel_index >= 4747) && (pixel_index <= 4793)) || ((pixel_index >= 4814) && (pixel_index <= 4831)) || ((pixel_index >= 4844) && (pixel_index <= 4889)) || ((pixel_index >= 4909) && (pixel_index <= 4927)) || ((pixel_index >= 4940) && (pixel_index <= 4985)) || ((pixel_index >= 5005) && (pixel_index <= 5023)) || ((pixel_index >= 5036) && (pixel_index <= 5081)) || ((pixel_index >= 5101) && (pixel_index <= 5119)) || ((pixel_index >= 5132) && (pixel_index <= 5177)) || ((pixel_index >= 5197) && (pixel_index <= 5215)) || ((pixel_index >= 5228) && (pixel_index <= 5273)) || ((pixel_index >= 5293) && (pixel_index <= 5311)) || ((pixel_index >= 5323) && (pixel_index <= 5369)) || pixel_index == 5381 || ((pixel_index >= 5389) && (pixel_index <= 5408)) || ((pixel_index >= 5419) && (pixel_index <= 5464)) || ((pixel_index >= 5477) && (pixel_index <= 5478)) || ((pixel_index >= 5486) && (pixel_index <= 5505)) || ((pixel_index >= 5514) && (pixel_index <= 5560)) || ((pixel_index >= 5573) && (pixel_index <= 5574)) || ((pixel_index >= 5582) && (pixel_index <= 5603)) || ((pixel_index >= 5608) && (pixel_index <= 5655)) || ((pixel_index >= 5669) && (pixel_index <= 5671)) || ((pixel_index >= 5678) && (pixel_index <= 5750)) || ((pixel_index >= 5765) && (pixel_index <= 5768)) || ((pixel_index >= 5774) && (pixel_index <= 5846)) || ((pixel_index >= 5861) && (pixel_index <= 5864)) || ((pixel_index >= 5871) && (pixel_index <= 5941)) || ((pixel_index >= 5957) && (pixel_index <= 5961)) || ((pixel_index >= 5967) && (pixel_index <= 6036)) || ((pixel_index >= 6053) && (pixel_index <= 6058)) || (pixel_index >= 6063) && (pixel_index <= 6131)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 5) begin
            if (((pixel_index >= 5) && (pixel_index <= 8)) || ((pixel_index >= 17) && (pixel_index <= 31)) || ((pixel_index >= 85) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 103)) || ((pixel_index >= 110) && (pixel_index <= 129)) || ((pixel_index >= 182) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 199)) || ((pixel_index >= 204) && (pixel_index <= 228)) || ((pixel_index >= 279) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 294)) || ((pixel_index >= 298) && (pixel_index <= 325)) || ((pixel_index >= 376) && (pixel_index <= 377)) || pixel_index == 389 || ((pixel_index >= 393) && (pixel_index <= 423)) || ((pixel_index >= 472) && (pixel_index <= 473)) || pixel_index == 485 || ((pixel_index >= 488) && (pixel_index <= 520)) || pixel_index == 569 || ((pixel_index >= 582) && (pixel_index <= 617)) || ((pixel_index >= 677) && (pixel_index <= 714)) || ((pixel_index >= 773) && (pixel_index <= 811)) || ((pixel_index >= 869) && (pixel_index <= 907)) || ((pixel_index >= 965) && (pixel_index <= 1004)) || ((pixel_index >= 1061) && (pixel_index <= 1100)) || ((pixel_index >= 1157) && (pixel_index <= 1197)) || ((pixel_index >= 1253) && (pixel_index <= 1293)) || ((pixel_index >= 1349) && (pixel_index <= 1390)) || ((pixel_index >= 1445) && (pixel_index <= 1486)) || ((pixel_index >= 1541) && (pixel_index <= 1583)) || ((pixel_index >= 1637) && (pixel_index <= 1656)) || ((pixel_index >= 1658) && (pixel_index <= 1679)) || ((pixel_index >= 1733) && (pixel_index <= 1749)) || ((pixel_index >= 1757) && (pixel_index <= 1775)) || ((pixel_index >= 1829) && (pixel_index <= 1844)) || ((pixel_index >= 1854) && (pixel_index <= 1871)) || ((pixel_index >= 1925) && (pixel_index <= 1939)) || ((pixel_index >= 1951) && (pixel_index <= 1967)) || ((pixel_index >= 2021) && (pixel_index <= 2035)) || ((pixel_index >= 2048) && (pixel_index <= 2064)) || ((pixel_index >= 2117) && (pixel_index <= 2131)) || ((pixel_index >= 2144) && (pixel_index <= 2160)) || ((pixel_index >= 2213) && (pixel_index <= 2226)) || ((pixel_index >= 2240) && (pixel_index <= 2256)) || ((pixel_index >= 2309) && (pixel_index <= 2322)) || ((pixel_index >= 2336) && (pixel_index <= 2352)) || ((pixel_index >= 2405) && (pixel_index <= 2419)) || ((pixel_index >= 2432) && (pixel_index <= 2448)) || ((pixel_index >= 2501) && (pixel_index <= 2515)) || ((pixel_index >= 2528) && (pixel_index <= 2544)) || ((pixel_index >= 2597) && (pixel_index <= 2611)) || ((pixel_index >= 2623) && (pixel_index <= 2639)) || ((pixel_index >= 2693) && (pixel_index <= 2708)) || ((pixel_index >= 2718) && (pixel_index <= 2735)) || ((pixel_index >= 2789) && (pixel_index <= 2806)) || ((pixel_index >= 2813) && (pixel_index <= 2831)) || ((pixel_index >= 2885) && (pixel_index <= 2927)) || ((pixel_index >= 2981) && (pixel_index <= 3023)) || ((pixel_index >= 3077) && (pixel_index <= 3118)) || ((pixel_index >= 3173) && (pixel_index <= 3214)) || ((pixel_index >= 3269) && (pixel_index <= 3310)) || ((pixel_index >= 3331) && (pixel_index <= 3335)) || ((pixel_index >= 3365) && (pixel_index <= 3405)) || ((pixel_index >= 3426) && (pixel_index <= 3433)) || ((pixel_index >= 3461) && (pixel_index <= 3501)) || ((pixel_index >= 3521) && (pixel_index <= 3529)) || ((pixel_index >= 3557) && (pixel_index <= 3597)) || ((pixel_index >= 3616) && (pixel_index <= 3626)) || ((pixel_index >= 3653) && (pixel_index <= 3693)) || ((pixel_index >= 3712) && (pixel_index <= 3722)) || ((pixel_index >= 3749) && (pixel_index <= 3789)) || ((pixel_index >= 3808) && (pixel_index <= 3818)) || ((pixel_index >= 3845) && (pixel_index <= 3885)) || ((pixel_index >= 3904) && (pixel_index <= 3914)) || ((pixel_index >= 3941) && (pixel_index <= 3981)) || ((pixel_index >= 4000) && (pixel_index <= 4010)) || ((pixel_index >= 4037) && (pixel_index <= 4077)) || ((pixel_index >= 4096) && (pixel_index <= 4106)) || ((pixel_index >= 4133) && (pixel_index <= 4173)) || ((pixel_index >= 4192) && (pixel_index <= 4201)) || ((pixel_index >= 4229) && (pixel_index <= 4269)) || ((pixel_index >= 4289) && (pixel_index <= 4296)) || ((pixel_index >= 4325) && (pixel_index <= 4366)) || ((pixel_index >= 4386) && (pixel_index <= 4391)) || ((pixel_index >= 4421) && (pixel_index <= 4462)) || ((pixel_index >= 4517) && (pixel_index <= 4558)) || ((pixel_index >= 4613) && (pixel_index <= 4654)) || ((pixel_index >= 4709) && (pixel_index <= 4751)) || ((pixel_index >= 4805) && (pixel_index <= 4847)) || ((pixel_index >= 4901) && (pixel_index <= 4944)) || ((pixel_index >= 4997) && (pixel_index <= 5040)) || ((pixel_index >= 5093) && (pixel_index <= 5137)) || ((pixel_index >= 5189) && (pixel_index <= 5234)) || ((pixel_index >= 5285) && (pixel_index <= 5330)) || ((pixel_index >= 5381) && (pixel_index <= 5427)) || ((pixel_index >= 5477) && (pixel_index <= 5524)) || pixel_index == 5561 || ((pixel_index >= 5573) && (pixel_index <= 5621)) || ((pixel_index >= 5655) && (pixel_index <= 5656)) || ((pixel_index >= 5670) && (pixel_index <= 5718)) || ((pixel_index >= 5750) && (pixel_index <= 5752)) || ((pixel_index >= 5767) && (pixel_index <= 5816)) || ((pixel_index >= 5845) && (pixel_index <= 5847)) || ((pixel_index >= 5863) && (pixel_index <= 5914)) || ((pixel_index >= 5939) && (pixel_index <= 5942)) || ((pixel_index >= 5960) && (pixel_index <= 6012)) || ((pixel_index >= 6033) && (pixel_index <= 6038)) || ((pixel_index >= 6057) && (pixel_index <= 6111)) || (pixel_index >= 6126) && (pixel_index <= 6133)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 6) begin
            if (((pixel_index >= 8) && (pixel_index <= 77)) || ((pixel_index >= 87) && (pixel_index <= 89)) || ((pixel_index >= 103) && (pixel_index <= 173)) || ((pixel_index >= 184) && (pixel_index <= 185)) || ((pixel_index >= 198) && (pixel_index <= 244)) || ((pixel_index >= 247) && (pixel_index <= 269)) || pixel_index == 281 || ((pixel_index >= 293) && (pixel_index <= 337)) || ((pixel_index >= 345) && (pixel_index <= 365)) || pixel_index == 377 || ((pixel_index >= 389) && (pixel_index <= 432)) || ((pixel_index >= 442) && (pixel_index <= 461)) || ((pixel_index >= 485) && (pixel_index <= 527)) || ((pixel_index >= 539) && (pixel_index <= 557)) || ((pixel_index >= 581) && (pixel_index <= 622)) || ((pixel_index >= 636) && (pixel_index <= 653)) || ((pixel_index >= 677) && (pixel_index <= 718)) || ((pixel_index >= 732) && (pixel_index <= 750)) || ((pixel_index >= 773) && (pixel_index <= 814)) || ((pixel_index >= 828) && (pixel_index <= 845)) || ((pixel_index >= 869) && (pixel_index <= 910)) || ((pixel_index >= 924) && (pixel_index <= 941)) || ((pixel_index >= 965) && (pixel_index <= 1006)) || ((pixel_index >= 1020) && (pixel_index <= 1037)) || ((pixel_index >= 1061) && (pixel_index <= 1102)) || ((pixel_index >= 1116) && (pixel_index <= 1133)) || ((pixel_index >= 1157) && (pixel_index <= 1199)) || ((pixel_index >= 1211) && (pixel_index <= 1229)) || ((pixel_index >= 1253) && (pixel_index <= 1296)) || ((pixel_index >= 1306) && (pixel_index <= 1325)) || ((pixel_index >= 1349) && (pixel_index <= 1393)) || ((pixel_index >= 1401) && (pixel_index <= 1420)) || ((pixel_index >= 1445) && (pixel_index <= 1492)) || ((pixel_index >= 1494) && (pixel_index <= 1516)) || ((pixel_index >= 1541) && (pixel_index <= 1612)) || ((pixel_index >= 1637) && (pixel_index <= 1707)) || ((pixel_index >= 1733) && (pixel_index <= 1803)) || ((pixel_index >= 1829) && (pixel_index <= 1898)) || ((pixel_index >= 1925) && (pixel_index <= 1994)) || ((pixel_index >= 2021) && (pixel_index <= 2089)) || ((pixel_index >= 2117) && (pixel_index <= 2184)) || ((pixel_index >= 2213) && (pixel_index <= 2280)) || ((pixel_index >= 2309) && (pixel_index <= 2375)) || ((pixel_index >= 2405) && (pixel_index <= 2470)) || ((pixel_index >= 2501) && (pixel_index <= 2565)) || ((pixel_index >= 2597) && (pixel_index <= 2660)) || ((pixel_index >= 2693) && (pixel_index <= 2754)) || ((pixel_index >= 2789) && (pixel_index <= 2848)) || ((pixel_index >= 2885) && (pixel_index <= 2942)) || ((pixel_index >= 2981) && (pixel_index <= 3013)) || ((pixel_index >= 3021) && (pixel_index <= 3035)) || ((pixel_index >= 3077) && (pixel_index <= 3105)) || ((pixel_index >= 3123) && (pixel_index <= 3126)) || ((pixel_index >= 3173) && (pixel_index <= 3199)) || ((pixel_index >= 3269) && (pixel_index <= 3292)) || ((pixel_index >= 3365) && (pixel_index <= 3387)) || ((pixel_index >= 3461) && (pixel_index <= 3481)) || ((pixel_index >= 3557) && (pixel_index <= 3576)) || ((pixel_index >= 3653) && (pixel_index <= 3671)) || ((pixel_index >= 3749) && (pixel_index <= 3766)) || ((pixel_index >= 3845) && (pixel_index <= 3861)) || ((pixel_index >= 3941) && (pixel_index <= 3956)) || ((pixel_index >= 4037) && (pixel_index <= 4052)) || ((pixel_index >= 4133) && (pixel_index <= 4147)) || ((pixel_index >= 4229) && (pixel_index <= 4242)) || ((pixel_index >= 4325) && (pixel_index <= 4338)) || ((pixel_index >= 4421) && (pixel_index <= 4434)) || ((pixel_index >= 4517) && (pixel_index <= 4529)) || ((pixel_index >= 4613) && (pixel_index <= 4625)) || ((pixel_index >= 4709) && (pixel_index <= 4721)) || ((pixel_index >= 4745) && (pixel_index <= 4746)) || ((pixel_index >= 4805) && (pixel_index <= 4816)) || ((pixel_index >= 4838) && (pixel_index <= 4844)) || ((pixel_index >= 4901) && (pixel_index <= 4912)) || ((pixel_index >= 4933) && (pixel_index <= 4941)) || ((pixel_index >= 4997) && (pixel_index <= 5008)) || ((pixel_index >= 5028) && (pixel_index <= 5038)) || ((pixel_index >= 5093) && (pixel_index <= 5104)) || ((pixel_index >= 5124) && (pixel_index <= 5135)) || ((pixel_index >= 5189) && (pixel_index <= 5200)) || ((pixel_index >= 5219) && (pixel_index <= 5231)) || ((pixel_index >= 5285) && (pixel_index <= 5296)) || ((pixel_index >= 5315) && (pixel_index <= 5327)) || ((pixel_index >= 5381) && (pixel_index <= 5392)) || ((pixel_index >= 5411) && (pixel_index <= 5423)) || ((pixel_index >= 5477) && (pixel_index <= 5488)) || ((pixel_index >= 5508) && (pixel_index <= 5519)) || ((pixel_index >= 5573) && (pixel_index <= 5584)) || ((pixel_index >= 5604) && (pixel_index <= 5614)) || ((pixel_index >= 5669) && (pixel_index <= 5680)) || ((pixel_index >= 5701) && (pixel_index <= 5709)) || ((pixel_index >= 5765) && (pixel_index <= 5776)) || ((pixel_index >= 5798) && (pixel_index <= 5804)) || pixel_index == 5849 || ((pixel_index >= 5862) && (pixel_index <= 5872)) || ((pixel_index >= 5944) && (pixel_index <= 5945)) || ((pixel_index >= 5959) && (pixel_index <= 5968)) || ((pixel_index >= 6040) && (pixel_index <= 6041)) || ((pixel_index >= 6056) && (pixel_index <= 6064)) || (pixel_index >= 6135) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 7) begin
            if (((pixel_index >= 6) && (pixel_index <= 88)) || ((pixel_index >= 101) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 377)) || ((pixel_index >= 389) && (pixel_index <= 399)) || ((pixel_index >= 411) && (pixel_index <= 473)) || ((pixel_index >= 485) && (pixel_index <= 492)) || ((pixel_index >= 511) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 586)) || ((pixel_index >= 609) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 680)) || ((pixel_index >= 707) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 775)) || ((pixel_index >= 804) && (pixel_index <= 857)) || pixel_index == 869 || ((pixel_index >= 902) && (pixel_index <= 953)) || ((pixel_index >= 999) && (pixel_index <= 1049)) || ((pixel_index >= 1096) && (pixel_index <= 1145)) || ((pixel_index >= 1193) && (pixel_index <= 1241)) || ((pixel_index >= 1290) && (pixel_index <= 1337)) || ((pixel_index >= 1386) && (pixel_index <= 1433)) || ((pixel_index >= 1483) && (pixel_index <= 1529)) || ((pixel_index >= 1580) && (pixel_index <= 1625)) || ((pixel_index >= 1676) && (pixel_index <= 1721)) || ((pixel_index >= 1773) && (pixel_index <= 1817)) || ((pixel_index >= 1869) && (pixel_index <= 1913)) || ((pixel_index >= 1966) && (pixel_index <= 2009)) || ((pixel_index >= 2062) && (pixel_index <= 2105)) || ((pixel_index >= 2159) && (pixel_index <= 2201)) || ((pixel_index >= 2229) && (pixel_index <= 2232)) || ((pixel_index >= 2255) && (pixel_index <= 2297)) || ((pixel_index >= 2323) && (pixel_index <= 2330)) || ((pixel_index >= 2351) && (pixel_index <= 2393)) || ((pixel_index >= 2418) && (pixel_index <= 2427)) || ((pixel_index >= 2447) && (pixel_index <= 2489)) || ((pixel_index >= 2514) && (pixel_index <= 2523)) || ((pixel_index >= 2543) && (pixel_index <= 2585)) || ((pixel_index >= 2609) && (pixel_index <= 2620)) || ((pixel_index >= 2640) && (pixel_index <= 2681)) || ((pixel_index >= 2705) && (pixel_index <= 2716)) || ((pixel_index >= 2736) && (pixel_index <= 2755)) || ((pixel_index >= 2763) && (pixel_index <= 2777)) || ((pixel_index >= 2801) && (pixel_index <= 2812)) || ((pixel_index >= 2832) && (pixel_index <= 2850)) || ((pixel_index >= 2860) && (pixel_index <= 2873)) || ((pixel_index >= 2897) && (pixel_index <= 2908)) || ((pixel_index >= 2928) && (pixel_index <= 2945)) || ((pixel_index >= 2957) && (pixel_index <= 2969)) || ((pixel_index >= 2993) && (pixel_index <= 3004)) || ((pixel_index >= 3024) && (pixel_index <= 3041)) || ((pixel_index >= 3054) && (pixel_index <= 3065)) || ((pixel_index >= 3089) && (pixel_index <= 3099)) || ((pixel_index >= 3120) && (pixel_index <= 3136)) || ((pixel_index >= 3150) && (pixel_index <= 3161)) || ((pixel_index >= 3186) && (pixel_index <= 3195)) || ((pixel_index >= 3215) && (pixel_index <= 3232)) || ((pixel_index >= 3246) && (pixel_index <= 3257)) || ((pixel_index >= 3283) && (pixel_index <= 3290)) || ((pixel_index >= 3312) && (pixel_index <= 3328)) || ((pixel_index >= 3342) && (pixel_index <= 3353)) || ((pixel_index >= 3380) && (pixel_index <= 3385)) || ((pixel_index >= 3408) && (pixel_index <= 3424)) || ((pixel_index >= 3438) && (pixel_index <= 3449)) || ((pixel_index >= 3504) && (pixel_index <= 3520)) || ((pixel_index >= 3534) && (pixel_index <= 3545)) || ((pixel_index >= 3600) && (pixel_index <= 3617)) || ((pixel_index >= 3630) && (pixel_index <= 3641)) || ((pixel_index >= 3696) && (pixel_index <= 3713)) || ((pixel_index >= 3725) && (pixel_index <= 3737)) || ((pixel_index >= 3792) && (pixel_index <= 3810)) || ((pixel_index >= 3820) && (pixel_index <= 3833)) || ((pixel_index >= 3888) && (pixel_index <= 3908)) || ((pixel_index >= 3915) && (pixel_index <= 3929)) || ((pixel_index >= 3985) && (pixel_index <= 4025)) || ((pixel_index >= 4081) && (pixel_index <= 4121)) || ((pixel_index >= 4178) && (pixel_index <= 4217)) || ((pixel_index >= 4274) && (pixel_index <= 4313)) || ((pixel_index >= 4370) && (pixel_index <= 4409)) || ((pixel_index >= 4467) && (pixel_index <= 4505)) || ((pixel_index >= 4563) && (pixel_index <= 4601)) || ((pixel_index >= 4660) && (pixel_index <= 4697)) || ((pixel_index >= 4757) && (pixel_index <= 4793)) || ((pixel_index >= 4853) && (pixel_index <= 4889)) || ((pixel_index >= 4950) && (pixel_index <= 4985)) || ((pixel_index >= 5047) && (pixel_index <= 5081)) || ((pixel_index >= 5145) && (pixel_index <= 5177)) || ((pixel_index >= 5242) && (pixel_index <= 5272)) || ((pixel_index >= 5339) && (pixel_index <= 5366)) || ((pixel_index >= 5437) && (pixel_index <= 5461)) || ((pixel_index >= 5534) && (pixel_index <= 5555)) || ((pixel_index >= 5633) && (pixel_index <= 5649)) || ((pixel_index >= 5733) && (pixel_index <= 5740)) || pixel_index == 5957 || pixel_index == 6041 || ((pixel_index >= 6053) && (pixel_index <= 6054)) || pixel_index == 6137) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 8) begin
            if (((pixel_index >= 67) && (pixel_index <= 89)) || ((pixel_index >= 135) && (pixel_index <= 139)) || ((pixel_index >= 164) && (pixel_index <= 185)) || ((pixel_index >= 229) && (pixel_index <= 237)) || ((pixel_index >= 260) && (pixel_index <= 281)) || ((pixel_index >= 324) && (pixel_index <= 333)) || ((pixel_index >= 356) && (pixel_index <= 377)) || ((pixel_index >= 420) && (pixel_index <= 430)) || ((pixel_index >= 452) && (pixel_index <= 473)) || ((pixel_index >= 515) && (pixel_index <= 527)) || ((pixel_index >= 548) && (pixel_index <= 569)) || ((pixel_index >= 611) && (pixel_index <= 623)) || ((pixel_index >= 644) && (pixel_index <= 665)) || ((pixel_index >= 707) && (pixel_index <= 719)) || ((pixel_index >= 740) && (pixel_index <= 761)) || ((pixel_index >= 803) && (pixel_index <= 815)) || ((pixel_index >= 836) && (pixel_index <= 857)) || ((pixel_index >= 899) && (pixel_index <= 910)) || ((pixel_index >= 932) && (pixel_index <= 953)) || ((pixel_index >= 996) && (pixel_index <= 1006)) || ((pixel_index >= 1028) && (pixel_index <= 1049)) || ((pixel_index >= 1092) && (pixel_index <= 1101)) || ((pixel_index >= 1124) && (pixel_index <= 1145)) || ((pixel_index >= 1189) && (pixel_index <= 1196)) || ((pixel_index >= 1219) && (pixel_index <= 1241)) || ((pixel_index >= 1288) && (pixel_index <= 1290)) || ((pixel_index >= 1315) && (pixel_index <= 1337)) || ((pixel_index >= 1411) && (pixel_index <= 1433)) || ((pixel_index >= 1506) && (pixel_index <= 1529)) || ((pixel_index >= 1602) && (pixel_index <= 1625)) || ((pixel_index >= 1697) && (pixel_index <= 1721)) || ((pixel_index >= 1793) && (pixel_index <= 1817)) || ((pixel_index >= 1888) && (pixel_index <= 1913)) || ((pixel_index >= 1984) && (pixel_index <= 2009)) || ((pixel_index >= 2079) && (pixel_index <= 2105)) || ((pixel_index >= 2174) && (pixel_index <= 2201)) || ((pixel_index >= 2270) && (pixel_index <= 2297)) || ((pixel_index >= 2365) && (pixel_index <= 2393)) || ((pixel_index >= 2460) && (pixel_index <= 2489)) || ((pixel_index >= 2555) && (pixel_index <= 2585)) || ((pixel_index >= 2650) && (pixel_index <= 2681)) || ((pixel_index >= 2744) && (pixel_index <= 2777)) || ((pixel_index >= 2839) && (pixel_index <= 2873)) || ((pixel_index >= 2932) && (pixel_index <= 2969)) || ((pixel_index >= 3026) && (pixel_index <= 3065)) || ((pixel_index >= 3118) && (pixel_index <= 3161)) || ((pixel_index >= 3211) && (pixel_index <= 3257)) || ((pixel_index >= 3305) && (pixel_index <= 3353)) || ((pixel_index >= 3400) && (pixel_index <= 3449)) || ((pixel_index >= 3494) && (pixel_index <= 3545)) || ((pixel_index >= 3589) && (pixel_index <= 3641)) || ((pixel_index >= 3684) && (pixel_index <= 3737)) || ((pixel_index >= 3779) && (pixel_index <= 3833)) || ((pixel_index >= 3874) && (pixel_index <= 3929)) || ((pixel_index >= 3969) && (pixel_index <= 4025)) || ((pixel_index >= 4064) && (pixel_index <= 4121)) || ((pixel_index >= 4159) && (pixel_index <= 4217)) || ((pixel_index >= 4255) && (pixel_index <= 4313)) || ((pixel_index >= 4350) && (pixel_index <= 4409)) || ((pixel_index >= 4446) && (pixel_index <= 4505)) || ((pixel_index >= 4541) && (pixel_index <= 4601)) || ((pixel_index >= 4637) && (pixel_index <= 4697)) || ((pixel_index >= 4732) && (pixel_index <= 4755)) || ((pixel_index >= 4759) && (pixel_index <= 4793)) || ((pixel_index >= 4828) && (pixel_index <= 4848)) || ((pixel_index >= 4857) && (pixel_index <= 4889)) || ((pixel_index >= 4924) && (pixel_index <= 4943)) || ((pixel_index >= 4954) && (pixel_index <= 4985)) || ((pixel_index >= 5020) && (pixel_index <= 5038)) || ((pixel_index >= 5051) && (pixel_index <= 5081)) || ((pixel_index >= 5115) && (pixel_index <= 5134)) || ((pixel_index >= 5148) && (pixel_index <= 5177)) || ((pixel_index >= 5211) && (pixel_index <= 5230)) || ((pixel_index >= 5244) && (pixel_index <= 5273)) || ((pixel_index >= 5307) && (pixel_index <= 5325)) || ((pixel_index >= 5340) && (pixel_index <= 5369)) || ((pixel_index >= 5403) && (pixel_index <= 5421)) || ((pixel_index >= 5436) && (pixel_index <= 5465)) || ((pixel_index >= 5499) && (pixel_index <= 5517)) || ((pixel_index >= 5532) && (pixel_index <= 5561)) || ((pixel_index >= 5595) && (pixel_index <= 5614)) || ((pixel_index >= 5628) && (pixel_index <= 5657)) || ((pixel_index >= 5691) && (pixel_index <= 5710)) || ((pixel_index >= 5724) && (pixel_index <= 5753)) || ((pixel_index >= 5787) && (pixel_index <= 5807)) || ((pixel_index >= 5819) && (pixel_index <= 5849)) || ((pixel_index >= 5883) && (pixel_index <= 5904)) || ((pixel_index >= 5914) && (pixel_index <= 5945)) || ((pixel_index >= 5980) && (pixel_index <= 6001)) || ((pixel_index >= 6008) && (pixel_index <= 6041)) || (pixel_index >= 6076) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 9) begin
            if (((pixel_index >= 445) && (pixel_index <= 446)) || ((pixel_index >= 538) && (pixel_index <= 545)) || ((pixel_index >= 633) && (pixel_index <= 642)) || ((pixel_index >= 729) && (pixel_index <= 739)) || ((pixel_index >= 824) && (pixel_index <= 835)) || ((pixel_index >= 920) && (pixel_index <= 931)) || ((pixel_index >= 1016) && (pixel_index <= 1027)) || ((pixel_index >= 1112) && (pixel_index <= 1123)) || ((pixel_index >= 1208) && (pixel_index <= 1219)) || ((pixel_index >= 1304) && (pixel_index <= 1315)) || ((pixel_index >= 1401) && (pixel_index <= 1410)) || ((pixel_index >= 1498) && (pixel_index <= 1505)) || ((pixel_index >= 1595) && (pixel_index <= 1600)) || ((pixel_index >= 2328) && (pixel_index <= 2336)) || ((pixel_index >= 2420) && (pixel_index <= 2436)) || ((pixel_index >= 2513) && (pixel_index <= 2534)) || ((pixel_index >= 2607) && (pixel_index <= 2632)) || pixel_index == 2681 || ((pixel_index >= 2702) && (pixel_index <= 2730)) || pixel_index == 2777 || ((pixel_index >= 2796) && (pixel_index <= 2827)) || ((pixel_index >= 2872) && (pixel_index <= 2873)) || ((pixel_index >= 2891) && (pixel_index <= 2925)) || ((pixel_index >= 2967) && (pixel_index <= 2969)) || ((pixel_index >= 2986) && (pixel_index <= 3022)) || ((pixel_index >= 3062) && (pixel_index <= 3065)) || ((pixel_index >= 3081) && (pixel_index <= 3119)) || ((pixel_index >= 3157) && (pixel_index <= 3161)) || ((pixel_index >= 3176) && (pixel_index <= 3216)) || ((pixel_index >= 3252) && (pixel_index <= 3257)) || ((pixel_index >= 3272) && (pixel_index <= 3313)) || ((pixel_index >= 3347) && (pixel_index <= 3353)) || ((pixel_index >= 3367) && (pixel_index <= 3410)) || ((pixel_index >= 3442) && (pixel_index <= 3449)) || ((pixel_index >= 3462) && (pixel_index <= 3508)) || ((pixel_index >= 3537) && (pixel_index <= 3545)) || ((pixel_index >= 3557) && (pixel_index <= 3606)) || ((pixel_index >= 3631) && (pixel_index <= 3641)) || ((pixel_index >= 3653) && (pixel_index <= 3704)) || ((pixel_index >= 3724) && (pixel_index <= 3737)) || ((pixel_index >= 3749) && (pixel_index <= 3803)) || ((pixel_index >= 3817) && (pixel_index <= 3833)) || ((pixel_index >= 3845) && (pixel_index <= 3929)) || ((pixel_index >= 3941) && (pixel_index <= 4025)) || ((pixel_index >= 4037) && (pixel_index <= 4121)) || ((pixel_index >= 4133) && (pixel_index <= 4217)) || ((pixel_index >= 4229) && (pixel_index <= 4313)) || ((pixel_index >= 4325) && (pixel_index <= 4351)) || ((pixel_index >= 4354) && (pixel_index <= 4409)) || ((pixel_index >= 4421) && (pixel_index <= 4444)) || ((pixel_index >= 4453) && (pixel_index <= 4505)) || ((pixel_index >= 4517) && (pixel_index <= 4539)) || ((pixel_index >= 4550) && (pixel_index <= 4601)) || ((pixel_index >= 4613) && (pixel_index <= 4634)) || ((pixel_index >= 4647) && (pixel_index <= 4697)) || ((pixel_index >= 4709) && (pixel_index <= 4729)) || ((pixel_index >= 4743) && (pixel_index <= 4793)) || ((pixel_index >= 4805) && (pixel_index <= 4825)) || ((pixel_index >= 4840) && (pixel_index <= 4889)) || ((pixel_index >= 4901) && (pixel_index <= 4921)) || ((pixel_index >= 4936) && (pixel_index <= 4985)) || ((pixel_index >= 4997) && (pixel_index <= 5017)) || ((pixel_index >= 5032) && (pixel_index <= 5081)) || ((pixel_index >= 5093) && (pixel_index <= 5113)) || ((pixel_index >= 5128) && (pixel_index <= 5177)) || ((pixel_index >= 5189) && (pixel_index <= 5209)) || ((pixel_index >= 5224) && (pixel_index <= 5273)) || ((pixel_index >= 5285) && (pixel_index <= 5305)) || ((pixel_index >= 5319) && (pixel_index <= 5369)) || ((pixel_index >= 5381) && (pixel_index <= 5402)) || ((pixel_index >= 5415) && (pixel_index <= 5465)) || ((pixel_index >= 5477) && (pixel_index <= 5499)) || ((pixel_index >= 5510) && (pixel_index <= 5561)) || ((pixel_index >= 5573) && (pixel_index <= 5596)) || ((pixel_index >= 5605) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5694)) || ((pixel_index >= 5699) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 6041)) || (pixel_index >= 6053) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 10) begin
            if (((pixel_index >= 595) && (pixel_index <= 597)) || ((pixel_index >= 685) && (pixel_index <= 699)) || ((pixel_index >= 778) && (pixel_index <= 798)) || ((pixel_index >= 872) && (pixel_index <= 896)) || ((pixel_index >= 967) && (pixel_index <= 994)) || ((pixel_index >= 1061) && (pixel_index <= 1091)) || ((pixel_index >= 1157) && (pixel_index <= 1189)) || ((pixel_index >= 1253) && (pixel_index <= 1286)) || ((pixel_index >= 1349) && (pixel_index <= 1383)) || ((pixel_index >= 1445) && (pixel_index <= 1480)) || ((pixel_index >= 1509) && (pixel_index <= 1513)) || ((pixel_index >= 1541) && (pixel_index <= 1576)) || ((pixel_index >= 1603) && (pixel_index <= 1611)) || ((pixel_index >= 1637) && (pixel_index <= 1673)) || ((pixel_index >= 1698) && (pixel_index <= 1707)) || ((pixel_index >= 1733) && (pixel_index <= 1770)) || ((pixel_index >= 1794) && (pixel_index <= 1804)) || ((pixel_index >= 1829) && (pixel_index <= 1867)) || ((pixel_index >= 1889) && (pixel_index <= 1901)) || ((pixel_index >= 1925) && (pixel_index <= 1963)) || ((pixel_index >= 1985) && (pixel_index <= 1997)) || ((pixel_index >= 2021) && (pixel_index <= 2060)) || ((pixel_index >= 2081) && (pixel_index <= 2093)) || ((pixel_index >= 2117) && (pixel_index <= 2156)) || ((pixel_index >= 2177) && (pixel_index <= 2189)) || ((pixel_index >= 2213) && (pixel_index <= 2252)) || ((pixel_index >= 2273) && (pixel_index <= 2285)) || ((pixel_index >= 2309) && (pixel_index <= 2349)) || ((pixel_index >= 2370) && (pixel_index <= 2380)) || ((pixel_index >= 2405) && (pixel_index <= 2445)) || ((pixel_index >= 2466) && (pixel_index <= 2476)) || ((pixel_index >= 2501) && (pixel_index <= 2542)) || ((pixel_index >= 2563) && (pixel_index <= 2571)) || ((pixel_index >= 2597) && (pixel_index <= 2638)) || ((pixel_index >= 2661) && (pixel_index <= 2665)) || ((pixel_index >= 2693) && (pixel_index <= 2734)) || ((pixel_index >= 2789) && (pixel_index <= 2830)) || ((pixel_index >= 2885) && (pixel_index <= 2926)) || ((pixel_index >= 2981) && (pixel_index <= 3022)) || ((pixel_index >= 3077) && (pixel_index <= 3118)) || ((pixel_index >= 3173) && (pixel_index <= 3214)) || ((pixel_index >= 3269) && (pixel_index <= 3311)) || ((pixel_index >= 3365) && (pixel_index <= 3379)) || ((pixel_index >= 3387) && (pixel_index <= 3407)) || ((pixel_index >= 3461) && (pixel_index <= 3474)) || ((pixel_index >= 3485) && (pixel_index <= 3503)) || ((pixel_index >= 3557) && (pixel_index <= 3569)) || ((pixel_index >= 3582) && (pixel_index <= 3599)) || ((pixel_index >= 3653) && (pixel_index <= 3664)) || ((pixel_index >= 3678) && (pixel_index <= 3695)) || ((pixel_index >= 3749) && (pixel_index <= 3760)) || ((pixel_index >= 3775) && (pixel_index <= 3792)) || ((pixel_index >= 3845) && (pixel_index <= 3856)) || ((pixel_index >= 3871) && (pixel_index <= 3888)) || ((pixel_index >= 3941) && (pixel_index <= 3952)) || ((pixel_index >= 3967) && (pixel_index <= 3984)) || ((pixel_index >= 4037) && (pixel_index <= 4048)) || ((pixel_index >= 4063) && (pixel_index <= 4081)) || ((pixel_index >= 4133) && (pixel_index <= 4144)) || ((pixel_index >= 4159) && (pixel_index <= 4177)) || ((pixel_index >= 4229) && (pixel_index <= 4240)) || ((pixel_index >= 4254) && (pixel_index <= 4274)) || ((pixel_index >= 4325) && (pixel_index <= 4337)) || ((pixel_index >= 4350) && (pixel_index <= 4370)) || ((pixel_index >= 4421) && (pixel_index <= 4433)) || ((pixel_index >= 4445) && (pixel_index <= 4467)) || ((pixel_index >= 4517) && (pixel_index <= 4530)) || ((pixel_index >= 4540) && (pixel_index <= 4564)) || ((pixel_index >= 4613) && (pixel_index <= 4628)) || ((pixel_index >= 4635) && (pixel_index <= 4661)) || ((pixel_index >= 4709) && (pixel_index <= 4758)) || ((pixel_index >= 4805) && (pixel_index <= 4854)) || ((pixel_index >= 4901) && (pixel_index <= 4952)) || ((pixel_index >= 4997) && (pixel_index <= 5049)) || ((pixel_index >= 5093) && (pixel_index <= 5146)) || pixel_index == 5177 || ((pixel_index >= 5189) && (pixel_index <= 5244)) || ((pixel_index >= 5272) && (pixel_index <= 5273)) || ((pixel_index >= 5285) && (pixel_index <= 5341)) || ((pixel_index >= 5366) && (pixel_index <= 5369)) || ((pixel_index >= 5381) && (pixel_index <= 5440)) || ((pixel_index >= 5459) && (pixel_index <= 5465)) || ((pixel_index >= 5477) && (pixel_index <= 5539)) || ((pixel_index >= 5552) && (pixel_index <= 5561)) || ((pixel_index >= 5573) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 6041)) || (pixel_index >= 6053) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 11) begin
            if (((pixel_index >= 5) && (pixel_index <= 40)) || ((pixel_index >= 101) && (pixel_index <= 137)) || ((pixel_index >= 197) && (pixel_index <= 234)) || ((pixel_index >= 293) && (pixel_index <= 331)) || ((pixel_index >= 389) && (pixel_index <= 428)) || ((pixel_index >= 485) && (pixel_index <= 524)) || ((pixel_index >= 581) && (pixel_index <= 621)) || ((pixel_index >= 677) && (pixel_index <= 717)) || ((pixel_index >= 773) && (pixel_index <= 814)) || ((pixel_index >= 869) && (pixel_index <= 910)) || ((pixel_index >= 965) && (pixel_index <= 1007)) || ((pixel_index >= 1061) && (pixel_index <= 1103)) || ((pixel_index >= 1157) && (pixel_index <= 1200)) || ((pixel_index >= 1253) && (pixel_index <= 1296)) || ((pixel_index >= 1349) && (pixel_index <= 1392)) || ((pixel_index >= 1445) && (pixel_index <= 1488)) || ((pixel_index >= 1541) && (pixel_index <= 1584)) || ((pixel_index >= 1637) && (pixel_index <= 1681)) || ((pixel_index >= 1733) && (pixel_index <= 1777)) || ((pixel_index >= 1829) && (pixel_index <= 1873)) || ((pixel_index >= 1925) && (pixel_index <= 1969)) || ((pixel_index >= 2021) && (pixel_index <= 2065)) || ((pixel_index >= 2117) && (pixel_index <= 2161)) || ((pixel_index >= 2213) && (pixel_index <= 2257)) || ((pixel_index >= 2279) && (pixel_index <= 2284)) || ((pixel_index >= 2309) && (pixel_index <= 2353)) || ((pixel_index >= 2374) && (pixel_index <= 2381)) || ((pixel_index >= 2405) && (pixel_index <= 2448)) || ((pixel_index >= 2469) && (pixel_index <= 2478)) || ((pixel_index >= 2501) && (pixel_index <= 2515)) || ((pixel_index >= 2519) && (pixel_index <= 2544)) || ((pixel_index >= 2564) && (pixel_index <= 2575)) || ((pixel_index >= 2597) && (pixel_index <= 2609)) || ((pixel_index >= 2617) && (pixel_index <= 2640)) || ((pixel_index >= 2660) && (pixel_index <= 2671)) || ((pixel_index >= 2693) && (pixel_index <= 2703)) || ((pixel_index >= 2715) && (pixel_index <= 2736)) || ((pixel_index >= 2756) && (pixel_index <= 2767)) || ((pixel_index >= 2789) && (pixel_index <= 2799)) || ((pixel_index >= 2811) && (pixel_index <= 2831)) || ((pixel_index >= 2852) && (pixel_index <= 2864)) || ((pixel_index >= 2885) && (pixel_index <= 2894)) || ((pixel_index >= 2908) && (pixel_index <= 2927)) || ((pixel_index >= 2948) && (pixel_index <= 2959)) || ((pixel_index >= 2981) && (pixel_index <= 2990)) || ((pixel_index >= 3004) && (pixel_index <= 3023)) || ((pixel_index >= 3044) && (pixel_index <= 3055)) || ((pixel_index >= 3077) && (pixel_index <= 3085)) || ((pixel_index >= 3101) && (pixel_index <= 3118)) || ((pixel_index >= 3140) && (pixel_index <= 3151)) || ((pixel_index >= 3173) && (pixel_index <= 3181)) || ((pixel_index >= 3197) && (pixel_index <= 3214)) || ((pixel_index >= 3237) && (pixel_index <= 3246)) || ((pixel_index >= 3269) && (pixel_index <= 3277)) || ((pixel_index >= 3293) && (pixel_index <= 3309)) || ((pixel_index >= 3334) && (pixel_index <= 3341)) || ((pixel_index >= 3365) && (pixel_index <= 3373)) || ((pixel_index >= 3388) && (pixel_index <= 3405)) || ((pixel_index >= 3432) && (pixel_index <= 3436)) || ((pixel_index >= 3461) && (pixel_index <= 3470)) || ((pixel_index >= 3484) && (pixel_index <= 3501)) || ((pixel_index >= 3557) && (pixel_index <= 3566)) || ((pixel_index >= 3580) && (pixel_index <= 3596)) || ((pixel_index >= 3653) && (pixel_index <= 3663)) || ((pixel_index >= 3675) && (pixel_index <= 3692)) || ((pixel_index >= 3749) && (pixel_index <= 3760)) || ((pixel_index >= 3770) && (pixel_index <= 3788)) || ((pixel_index >= 3845) && (pixel_index <= 3857)) || ((pixel_index >= 3865) && (pixel_index <= 3884)) || ((pixel_index >= 3941) && (pixel_index <= 3980)) || ((pixel_index >= 4037) && (pixel_index <= 4076)) || ((pixel_index >= 4133) && (pixel_index <= 4172)) || ((pixel_index >= 4229) && (pixel_index <= 4268)) || ((pixel_index >= 4325) && (pixel_index <= 4364)) || ((pixel_index >= 4421) && (pixel_index <= 4460)) || ((pixel_index >= 4517) && (pixel_index <= 4556)) || ((pixel_index >= 4613) && (pixel_index <= 4652)) || ((pixel_index >= 4709) && (pixel_index <= 4748)) || ((pixel_index >= 4805) && (pixel_index <= 4845)) || ((pixel_index >= 4901) && (pixel_index <= 4941)) || ((pixel_index >= 4997) && (pixel_index <= 5037)) || ((pixel_index >= 5093) && (pixel_index <= 5133)) || ((pixel_index >= 5189) && (pixel_index <= 5230)) || ((pixel_index >= 5285) && (pixel_index <= 5326)) || ((pixel_index >= 5381) && (pixel_index <= 5423)) || ((pixel_index >= 5477) && (pixel_index <= 5519)) || ((pixel_index >= 5573) && (pixel_index <= 5616)) || ((pixel_index >= 5669) && (pixel_index <= 5713)) || ((pixel_index >= 5765) && (pixel_index <= 5809)) || ((pixel_index >= 5861) && (pixel_index <= 5906)) || ((pixel_index >= 5957) && (pixel_index <= 6003)) || (pixel_index >= 6053) && (pixel_index <= 6100)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 12) begin
            if (((pixel_index >= 5) && (pixel_index <= 46)) || ((pixel_index >= 101) && (pixel_index <= 142)) || ((pixel_index >= 197) && (pixel_index <= 238)) || ((pixel_index >= 293) && (pixel_index <= 335)) || ((pixel_index >= 389) && (pixel_index <= 431)) || ((pixel_index >= 485) && (pixel_index <= 527)) || ((pixel_index >= 581) && (pixel_index <= 623)) || ((pixel_index >= 677) && (pixel_index <= 719)) || ((pixel_index >= 773) && (pixel_index <= 815)) || ((pixel_index >= 869) && (pixel_index <= 911)) || ((pixel_index >= 965) && (pixel_index <= 1007)) || ((pixel_index >= 1061) && (pixel_index <= 1103)) || ((pixel_index >= 1157) && (pixel_index <= 1199)) || ((pixel_index >= 1253) && (pixel_index <= 1295)) || ((pixel_index >= 1349) && (pixel_index <= 1391)) || ((pixel_index >= 1445) && (pixel_index <= 1487)) || ((pixel_index >= 1541) && (pixel_index <= 1583)) || ((pixel_index >= 1637) && (pixel_index <= 1679)) || ((pixel_index >= 1733) && (pixel_index <= 1775)) || ((pixel_index >= 1829) && (pixel_index <= 1871)) || ((pixel_index >= 1925) && (pixel_index <= 1967)) || ((pixel_index >= 2021) && (pixel_index <= 2063)) || ((pixel_index >= 2117) && (pixel_index <= 2159)) || ((pixel_index >= 2213) && (pixel_index <= 2255)) || ((pixel_index >= 2309) && (pixel_index <= 2322)) || ((pixel_index >= 2328) && (pixel_index <= 2351)) || ((pixel_index >= 2405) && (pixel_index <= 2416)) || ((pixel_index >= 2426) && (pixel_index <= 2447)) || ((pixel_index >= 2473) && (pixel_index <= 2475)) || ((pixel_index >= 2501) && (pixel_index <= 2511)) || ((pixel_index >= 2523) && (pixel_index <= 2543)) || ((pixel_index >= 2567) && (pixel_index <= 2573)) || ((pixel_index >= 2597) && (pixel_index <= 2606)) || ((pixel_index >= 2619) && (pixel_index <= 2639)) || ((pixel_index >= 2661) && (pixel_index <= 2670)) || ((pixel_index >= 2693) && (pixel_index <= 2702)) || ((pixel_index >= 2716) && (pixel_index <= 2735)) || ((pixel_index >= 2757) && (pixel_index <= 2767)) || ((pixel_index >= 2789) && (pixel_index <= 2797)) || ((pixel_index >= 2812) && (pixel_index <= 2831)) || ((pixel_index >= 2852) && (pixel_index <= 2863)) || ((pixel_index >= 2885) && (pixel_index <= 2893)) || ((pixel_index >= 2908) && (pixel_index <= 2927)) || ((pixel_index >= 2948) && (pixel_index <= 2960)) || ((pixel_index >= 2981) && (pixel_index <= 2989)) || ((pixel_index >= 3005) && (pixel_index <= 3023)) || ((pixel_index >= 3044) && (pixel_index <= 3056)) || ((pixel_index >= 3077) && (pixel_index <= 3085)) || ((pixel_index >= 3100) && (pixel_index <= 3118)) || ((pixel_index >= 3140) && (pixel_index <= 3152)) || ((pixel_index >= 3173) && (pixel_index <= 3181)) || ((pixel_index >= 3196) && (pixel_index <= 3214)) || ((pixel_index >= 3236) && (pixel_index <= 3248)) || ((pixel_index >= 3269) && (pixel_index <= 3278)) || ((pixel_index >= 3292) && (pixel_index <= 3310)) || ((pixel_index >= 3332) && (pixel_index <= 3343)) || ((pixel_index >= 3365) && (pixel_index <= 3374)) || ((pixel_index >= 3387) && (pixel_index <= 3406)) || ((pixel_index >= 3429) && (pixel_index <= 3439)) || ((pixel_index >= 3461) && (pixel_index <= 3471)) || ((pixel_index >= 3483) && (pixel_index <= 3502)) || ((pixel_index >= 3526) && (pixel_index <= 3534)) || ((pixel_index >= 3557) && (pixel_index <= 3568)) || ((pixel_index >= 3578) && (pixel_index <= 3598)) || ((pixel_index >= 3623) && (pixel_index <= 3628)) || ((pixel_index >= 3653) && (pixel_index <= 3666)) || ((pixel_index >= 3672) && (pixel_index <= 3694)) || ((pixel_index >= 3749) && (pixel_index <= 3790)) || ((pixel_index >= 3845) && (pixel_index <= 3886)) || ((pixel_index >= 3941) && (pixel_index <= 3982)) || ((pixel_index >= 4037) && (pixel_index <= 4078)) || ((pixel_index >= 4133) && (pixel_index <= 4174)) || ((pixel_index >= 4229) && (pixel_index <= 4270)) || ((pixel_index >= 4325) && (pixel_index <= 4366)) || ((pixel_index >= 4421) && (pixel_index <= 4462)) || ((pixel_index >= 4517) && (pixel_index <= 4558)) || ((pixel_index >= 4613) && (pixel_index <= 4654)) || ((pixel_index >= 4709) && (pixel_index <= 4750)) || ((pixel_index >= 4805) && (pixel_index <= 4846)) || ((pixel_index >= 4901) && (pixel_index <= 4942)) || ((pixel_index >= 4997) && (pixel_index <= 5038)) || ((pixel_index >= 5093) && (pixel_index <= 5134)) || ((pixel_index >= 5189) && (pixel_index <= 5230)) || ((pixel_index >= 5285) && (pixel_index <= 5326)) || ((pixel_index >= 5381) && (pixel_index <= 5422)) || ((pixel_index >= 5477) && (pixel_index <= 5518)) || ((pixel_index >= 5573) && (pixel_index <= 5614)) || ((pixel_index >= 5669) && (pixel_index <= 5711)) || ((pixel_index >= 5765) && (pixel_index <= 5807)) || ((pixel_index >= 5861) && (pixel_index <= 5903)) || ((pixel_index >= 5957) && (pixel_index <= 5999)) || (pixel_index >= 6053) && (pixel_index <= 6095)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 13) begin
            if (((pixel_index >= 5) && (pixel_index <= 38)) || ((pixel_index >= 101) && (pixel_index <= 134)) || ((pixel_index >= 197) && (pixel_index <= 230)) || ((pixel_index >= 293) && (pixel_index <= 326)) || ((pixel_index >= 389) && (pixel_index <= 422)) || ((pixel_index >= 485) && (pixel_index <= 518)) || ((pixel_index >= 581) && (pixel_index <= 614)) || ((pixel_index >= 677) && (pixel_index <= 710)) || ((pixel_index >= 773) && (pixel_index <= 806)) || ((pixel_index >= 869) && (pixel_index <= 902)) || ((pixel_index >= 965) && (pixel_index <= 998)) || ((pixel_index >= 1061) && (pixel_index <= 1094)) || ((pixel_index >= 1157) && (pixel_index <= 1190)) || ((pixel_index >= 1253) && (pixel_index <= 1286)) || ((pixel_index >= 1349) && (pixel_index <= 1382)) || ((pixel_index >= 1445) && (pixel_index <= 1478)) || ((pixel_index >= 1541) && (pixel_index <= 1574)) || ((pixel_index >= 1637) && (pixel_index <= 1670)) || ((pixel_index >= 1733) && (pixel_index <= 1766)) || ((pixel_index >= 1829) && (pixel_index <= 1862)) || ((pixel_index >= 1925) && (pixel_index <= 1958)) || ((pixel_index >= 2021) && (pixel_index <= 2054)) || ((pixel_index >= 2117) && (pixel_index <= 2150)) || ((pixel_index >= 2213) && (pixel_index <= 2246)) || ((pixel_index >= 2309) && (pixel_index <= 2314)) || ((pixel_index >= 2319) && (pixel_index <= 2342)) || ((pixel_index >= 2405) && (pixel_index <= 2408)) || ((pixel_index >= 2417) && (pixel_index <= 2438)) || ((pixel_index >= 2464) && (pixel_index <= 2467)) || ((pixel_index >= 2501) && (pixel_index <= 2503)) || ((pixel_index >= 2514) && (pixel_index <= 2534)) || ((pixel_index >= 2558) && (pixel_index <= 2565)) || ((pixel_index >= 2597) && (pixel_index <= 2598)) || ((pixel_index >= 2611) && (pixel_index <= 2630)) || ((pixel_index >= 2653) && (pixel_index <= 2662)) || ((pixel_index >= 2693) && (pixel_index <= 2694)) || ((pixel_index >= 2708) && (pixel_index <= 2726)) || ((pixel_index >= 2748) && (pixel_index <= 2759)) || pixel_index == 2789 || ((pixel_index >= 2804) && (pixel_index <= 2822)) || ((pixel_index >= 2843) && (pixel_index <= 2856)) || pixel_index == 2885 || ((pixel_index >= 2900) && (pixel_index <= 2918)) || ((pixel_index >= 2939) && (pixel_index <= 2958)) || pixel_index == 2981 || ((pixel_index >= 2996) && (pixel_index <= 3014)) || ((pixel_index >= 3031) && (pixel_index <= 3056)) || pixel_index == 3077 || ((pixel_index >= 3092) && (pixel_index <= 3110)) || ((pixel_index >= 3125) && (pixel_index <= 3152)) || pixel_index == 3173 || ((pixel_index >= 3188) && (pixel_index <= 3206)) || ((pixel_index >= 3223) && (pixel_index <= 3247)) || ((pixel_index >= 3269) && (pixel_index <= 3270)) || ((pixel_index >= 3284) && (pixel_index <= 3302)) || ((pixel_index >= 3323) && (pixel_index <= 3336)) || ((pixel_index >= 3338) && (pixel_index <= 3342)) || ((pixel_index >= 3365) && (pixel_index <= 3366)) || ((pixel_index >= 3379) && (pixel_index <= 3398)) || ((pixel_index >= 3420) && (pixel_index <= 3431)) || ((pixel_index >= 3461) && (pixel_index <= 3463)) || ((pixel_index >= 3474) && (pixel_index <= 3494)) || ((pixel_index >= 3517) && (pixel_index <= 3526)) || ((pixel_index >= 3557) && (pixel_index <= 3560)) || ((pixel_index >= 3569) && (pixel_index <= 3590)) || ((pixel_index >= 3614) && (pixel_index <= 3620)) || ((pixel_index >= 3653) && (pixel_index <= 3658)) || ((pixel_index >= 3663) && (pixel_index <= 3686)) || ((pixel_index >= 3749) && (pixel_index <= 3782)) || ((pixel_index >= 3845) && (pixel_index <= 3878)) || ((pixel_index >= 3941) && (pixel_index <= 3974)) || ((pixel_index >= 4037) && (pixel_index <= 4070)) || ((pixel_index >= 4133) && (pixel_index <= 4166)) || ((pixel_index >= 4229) && (pixel_index <= 4262)) || ((pixel_index >= 4325) && (pixel_index <= 4358)) || ((pixel_index >= 4421) && (pixel_index <= 4454)) || ((pixel_index >= 4517) && (pixel_index <= 4550)) || ((pixel_index >= 4613) && (pixel_index <= 4646)) || ((pixel_index >= 4709) && (pixel_index <= 4742)) || ((pixel_index >= 4805) && (pixel_index <= 4838)) || ((pixel_index >= 4901) && (pixel_index <= 4934)) || ((pixel_index >= 4997) && (pixel_index <= 5030)) || ((pixel_index >= 5093) && (pixel_index <= 5126)) || ((pixel_index >= 5189) && (pixel_index <= 5222)) || ((pixel_index >= 5285) && (pixel_index <= 5318)) || ((pixel_index >= 5381) && (pixel_index <= 5414)) || ((pixel_index >= 5477) && (pixel_index <= 5510)) || ((pixel_index >= 5573) && (pixel_index <= 5606)) || ((pixel_index >= 5669) && (pixel_index <= 5702)) || ((pixel_index >= 5765) && (pixel_index <= 5798)) || ((pixel_index >= 5861) && (pixel_index <= 5894)) || ((pixel_index >= 5957) && (pixel_index <= 5990)) || (pixel_index >= 6053) && (pixel_index <= 6086)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 14) begin
            if (((pixel_index >= 5) && (pixel_index <= 29)) || ((pixel_index >= 101) && (pixel_index <= 125)) || ((pixel_index >= 197) && (pixel_index <= 221)) || ((pixel_index >= 293) && (pixel_index <= 317)) || ((pixel_index >= 389) && (pixel_index <= 413)) || ((pixel_index >= 485) && (pixel_index <= 509)) || ((pixel_index >= 581) && (pixel_index <= 605)) || ((pixel_index >= 677) && (pixel_index <= 701)) || ((pixel_index >= 773) && (pixel_index <= 797)) || ((pixel_index >= 869) && (pixel_index <= 893)) || ((pixel_index >= 965) && (pixel_index <= 989)) || ((pixel_index >= 1061) && (pixel_index <= 1085)) || ((pixel_index >= 1157) && (pixel_index <= 1181)) || ((pixel_index >= 1253) && (pixel_index <= 1277)) || ((pixel_index >= 1349) && (pixel_index <= 1373)) || ((pixel_index >= 1445) && (pixel_index <= 1469)) || ((pixel_index >= 1541) && (pixel_index <= 1565)) || ((pixel_index >= 1637) && (pixel_index <= 1661)) || ((pixel_index >= 1733) && (pixel_index <= 1757)) || ((pixel_index >= 1829) && (pixel_index <= 1853)) || ((pixel_index >= 1925) && (pixel_index <= 1949)) || ((pixel_index >= 2021) && (pixel_index <= 2045)) || ((pixel_index >= 2117) && (pixel_index <= 2141)) || ((pixel_index >= 2168) && (pixel_index <= 2170)) || ((pixel_index >= 2213) && (pixel_index <= 2237)) || ((pixel_index >= 2260) && (pixel_index <= 2269)) || ((pixel_index >= 2310) && (pixel_index <= 2333)) || ((pixel_index >= 2354) && (pixel_index <= 2367)) || ((pixel_index >= 2408) && (pixel_index <= 2429)) || ((pixel_index >= 2449) && (pixel_index <= 2463)) || ((pixel_index >= 2505) && (pixel_index <= 2525)) || ((pixel_index >= 2544) && (pixel_index <= 2560)) || ((pixel_index >= 2602) && (pixel_index <= 2621)) || ((pixel_index >= 2640) && (pixel_index <= 2656)) || ((pixel_index >= 2698) && (pixel_index <= 2717)) || ((pixel_index >= 2736) && (pixel_index <= 2753)) || ((pixel_index >= 2795) && (pixel_index <= 2813)) || ((pixel_index >= 2832) && (pixel_index <= 2849)) || ((pixel_index >= 2891) && (pixel_index <= 2909)) || ((pixel_index >= 2929) && (pixel_index <= 2945)) || ((pixel_index >= 2957) && (pixel_index <= 2959)) || ((pixel_index >= 2987) && (pixel_index <= 3005)) || ((pixel_index >= 3025) && (pixel_index <= 3044)) || ((pixel_index >= 3046) && (pixel_index <= 3056)) || ((pixel_index >= 3083) && (pixel_index <= 3101)) || ((pixel_index >= 3122) && (pixel_index <= 3154)) || ((pixel_index >= 3179) && (pixel_index <= 3197)) || ((pixel_index >= 3203) && (pixel_index <= 3215)) || ((pixel_index >= 3218) && (pixel_index <= 3251)) || ((pixel_index >= 3274) && (pixel_index <= 3293)) || ((pixel_index >= 3299) && (pixel_index <= 3347)) || ((pixel_index >= 3370) && (pixel_index <= 3389)) || ((pixel_index >= 3399) && (pixel_index <= 3400)) || ((pixel_index >= 3414) && (pixel_index <= 3443)) || ((pixel_index >= 3465) && (pixel_index <= 3485)) || ((pixel_index >= 3511) && (pixel_index <= 3539)) || ((pixel_index >= 3560) && (pixel_index <= 3581)) || ((pixel_index >= 3608) && (pixel_index <= 3620)) || ((pixel_index >= 3623) && (pixel_index <= 3633)) || ((pixel_index >= 3654) && (pixel_index <= 3677)) || ((pixel_index >= 3705) && (pixel_index <= 3715)) || ((pixel_index >= 3723) && (pixel_index <= 3728)) || ((pixel_index >= 3749) && (pixel_index <= 3773)) || ((pixel_index >= 3802) && (pixel_index <= 3810)) || pixel_index == 3823 || ((pixel_index >= 3845) && (pixel_index <= 3869)) || ((pixel_index >= 3941) && (pixel_index <= 3965)) || ((pixel_index >= 4037) && (pixel_index <= 4061)) || ((pixel_index >= 4133) && (pixel_index <= 4157)) || ((pixel_index >= 4229) && (pixel_index <= 4253)) || ((pixel_index >= 4325) && (pixel_index <= 4349)) || ((pixel_index >= 4421) && (pixel_index <= 4445)) || ((pixel_index >= 4517) && (pixel_index <= 4541)) || ((pixel_index >= 4613) && (pixel_index <= 4637)) || ((pixel_index >= 4709) && (pixel_index <= 4733)) || ((pixel_index >= 4805) && (pixel_index <= 4829)) || ((pixel_index >= 4901) && (pixel_index <= 4925)) || ((pixel_index >= 4997) && (pixel_index <= 5021)) || ((pixel_index >= 5093) && (pixel_index <= 5117)) || ((pixel_index >= 5189) && (pixel_index <= 5213)) || ((pixel_index >= 5285) && (pixel_index <= 5309)) || ((pixel_index >= 5381) && (pixel_index <= 5405)) || ((pixel_index >= 5477) && (pixel_index <= 5501)) || ((pixel_index >= 5573) && (pixel_index <= 5597)) || ((pixel_index >= 5669) && (pixel_index <= 5693)) || ((pixel_index >= 5765) && (pixel_index <= 5789)) || ((pixel_index >= 5861) && (pixel_index <= 5885)) || ((pixel_index >= 5957) && (pixel_index <= 5981)) || (pixel_index >= 6053) && (pixel_index <= 6077)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 15) begin
            if (((pixel_index >= 5) && (pixel_index <= 25)) || ((pixel_index >= 101) && (pixel_index <= 121)) || ((pixel_index >= 197) && (pixel_index <= 217)) || ((pixel_index >= 293) && (pixel_index <= 313)) || ((pixel_index >= 389) && (pixel_index <= 409)) || ((pixel_index >= 485) && (pixel_index <= 505)) || ((pixel_index >= 581) && (pixel_index <= 601)) || ((pixel_index >= 677) && (pixel_index <= 697)) || ((pixel_index >= 773) && (pixel_index <= 793)) || ((pixel_index >= 869) && (pixel_index <= 889)) || ((pixel_index >= 965) && (pixel_index <= 985)) || ((pixel_index >= 1061) && (pixel_index <= 1081)) || ((pixel_index >= 1157) && (pixel_index <= 1177)) || ((pixel_index >= 1253) && (pixel_index <= 1273)) || ((pixel_index >= 1349) && (pixel_index <= 1369)) || ((pixel_index >= 1445) && (pixel_index <= 1465)) || ((pixel_index >= 1541) && (pixel_index <= 1561)) || ((pixel_index >= 1637) && (pixel_index <= 1657)) || ((pixel_index >= 1733) && (pixel_index <= 1753)) || ((pixel_index >= 1783) && (pixel_index <= 1786)) || ((pixel_index >= 1829) && (pixel_index <= 1849)) || ((pixel_index >= 1877) && (pixel_index <= 1883)) || ((pixel_index >= 1925) && (pixel_index <= 1945)) || ((pixel_index >= 1973) && (pixel_index <= 1981)) || ((pixel_index >= 2021) && (pixel_index <= 2041)) || ((pixel_index >= 2063) && (pixel_index <= 2064)) || ((pixel_index >= 2067) && (pixel_index <= 2074)) || ((pixel_index >= 2077) && (pixel_index <= 2078)) || ((pixel_index >= 2117) && (pixel_index <= 2137)) || ((pixel_index >= 2159) && (pixel_index <= 2170)) || ((pixel_index >= 2213) && (pixel_index <= 2233)) || ((pixel_index >= 2255) && (pixel_index <= 2270)) || ((pixel_index >= 2309) && (pixel_index <= 2329)) || ((pixel_index >= 2351) && (pixel_index <= 2367)) || ((pixel_index >= 2405) && (pixel_index <= 2425)) || ((pixel_index >= 2449) && (pixel_index <= 2464)) || ((pixel_index >= 2501) && (pixel_index <= 2521)) || ((pixel_index >= 2548) && (pixel_index <= 2562)) || ((pixel_index >= 2598) && (pixel_index <= 2617)) || ((pixel_index >= 2647) && (pixel_index <= 2658)) || ((pixel_index >= 2695) && (pixel_index <= 2713)) || ((pixel_index >= 2743) && (pixel_index <= 2754)) || ((pixel_index >= 2791) && (pixel_index <= 2809)) || ((pixel_index >= 2839) && (pixel_index <= 2848)) || ((pixel_index >= 2887) && (pixel_index <= 2905)) || ((pixel_index >= 2935) && (pixel_index <= 2940)) || ((pixel_index >= 2943) && (pixel_index <= 2944)) || ((pixel_index >= 2983) && (pixel_index <= 3001)) || ((pixel_index >= 3030) && (pixel_index <= 3036)) || ((pixel_index >= 3038) && (pixel_index <= 3040)) || ((pixel_index >= 3079) && (pixel_index <= 3097)) || ((pixel_index >= 3127) && (pixel_index <= 3136)) || ((pixel_index >= 3175) && (pixel_index <= 3193)) || ((pixel_index >= 3222) && (pixel_index <= 3232)) || ((pixel_index >= 3271) && (pixel_index <= 3289)) || ((pixel_index >= 3318) && (pixel_index <= 3319)) || ((pixel_index >= 3321) && (pixel_index <= 3332)) || ((pixel_index >= 3366) && (pixel_index <= 3385)) || ((pixel_index >= 3413) && (pixel_index <= 3415)) || ((pixel_index >= 3417) && (pixel_index <= 3431)) || ((pixel_index >= 3437) && (pixel_index <= 3438)) || ((pixel_index >= 3461) && (pixel_index <= 3481)) || ((pixel_index >= 3509) && (pixel_index <= 3510)) || ((pixel_index >= 3513) && (pixel_index <= 3537)) || ((pixel_index >= 3557) && (pixel_index <= 3577)) || ((pixel_index >= 3583) && (pixel_index <= 3589)) || ((pixel_index >= 3604) && (pixel_index <= 3605)) || ((pixel_index >= 3607) && (pixel_index <= 3634)) || ((pixel_index >= 3653) && (pixel_index <= 3673)) || ((pixel_index >= 3679) && (pixel_index <= 3731)) || ((pixel_index >= 3749) && (pixel_index <= 3769)) || ((pixel_index >= 3778) && (pixel_index <= 3828)) || ((pixel_index >= 3845) && (pixel_index <= 3865)) || pixel_index == 3876 || ((pixel_index >= 3880) && (pixel_index <= 3883)) || ((pixel_index >= 3892) && (pixel_index <= 3925)) || ((pixel_index >= 3941) && (pixel_index <= 3961)) || ((pixel_index >= 3978) && (pixel_index <= 3979)) || ((pixel_index >= 3990) && (pixel_index <= 4021)) || ((pixel_index >= 4037) && (pixel_index <= 4057)) || pixel_index == 4075 || ((pixel_index >= 4085) && (pixel_index <= 4117)) || ((pixel_index >= 4133) && (pixel_index <= 4153)) || pixel_index == 4172 || pixel_index == 4183 || ((pixel_index >= 4185) && (pixel_index <= 4194)) || ((pixel_index >= 4200) && (pixel_index <= 4212)) || ((pixel_index >= 4229) && (pixel_index <= 4249)) || ((pixel_index >= 4285) && (pixel_index <= 4288)) || ((pixel_index >= 4301) && (pixel_index <= 4306)) || ((pixel_index >= 4325) && (pixel_index <= 4345)) || ((pixel_index >= 4382) && (pixel_index <= 4384)) || ((pixel_index >= 4399) && (pixel_index <= 4401)) || ((pixel_index >= 4421) && (pixel_index <= 4441)) || ((pixel_index >= 4479) && (pixel_index <= 4480)) || ((pixel_index >= 4517) && (pixel_index <= 4537)) || ((pixel_index >= 4613) && (pixel_index <= 4633)) || ((pixel_index >= 4709) && (pixel_index <= 4729)) || ((pixel_index >= 4805) && (pixel_index <= 4825)) || ((pixel_index >= 4901) && (pixel_index <= 4921)) || ((pixel_index >= 4997) && (pixel_index <= 5017)) || ((pixel_index >= 5093) && (pixel_index <= 5113)) || ((pixel_index >= 5189) && (pixel_index <= 5209)) || ((pixel_index >= 5285) && (pixel_index <= 5305)) || ((pixel_index >= 5381) && (pixel_index <= 5401)) || ((pixel_index >= 5477) && (pixel_index <= 5497)) || ((pixel_index >= 5573) && (pixel_index <= 5593)) || ((pixel_index >= 5669) && (pixel_index <= 5689)) || ((pixel_index >= 5765) && (pixel_index <= 5785)) || ((pixel_index >= 5861) && (pixel_index <= 5881)) || ((pixel_index >= 5957) && (pixel_index <= 5977)) || (pixel_index >= 6053) && (pixel_index <= 6073)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 16) begin
            if (((pixel_index >= 5) && (pixel_index <= 22)) || ((pixel_index >= 101) && (pixel_index <= 118)) || ((pixel_index >= 197) && (pixel_index <= 214)) || ((pixel_index >= 293) && (pixel_index <= 310)) || ((pixel_index >= 389) && (pixel_index <= 406)) || ((pixel_index >= 485) && (pixel_index <= 502)) || ((pixel_index >= 581) && (pixel_index <= 598)) || ((pixel_index >= 677) && (pixel_index <= 694)) || ((pixel_index >= 773) && (pixel_index <= 790)) || ((pixel_index >= 869) && (pixel_index <= 886)) || ((pixel_index >= 965) && (pixel_index <= 982)) || ((pixel_index >= 1061) && (pixel_index <= 1078)) || ((pixel_index >= 1157) && (pixel_index <= 1174)) || ((pixel_index >= 1253) && (pixel_index <= 1270)) || ((pixel_index >= 1349) && (pixel_index <= 1366)) || ((pixel_index >= 1445) && (pixel_index <= 1462)) || ((pixel_index >= 1541) && (pixel_index <= 1558)) || ((pixel_index >= 1637) && (pixel_index <= 1654)) || ((pixel_index >= 1733) && (pixel_index <= 1750)) || ((pixel_index >= 1829) && (pixel_index <= 1846)) || ((pixel_index >= 1925) && (pixel_index <= 1942)) || ((pixel_index >= 2021) && (pixel_index <= 2038)) || ((pixel_index >= 2069) && (pixel_index <= 2072)) || ((pixel_index >= 2117) && (pixel_index <= 2134)) || ((pixel_index >= 2164) && (pixel_index <= 2170)) || ((pixel_index >= 2213) && (pixel_index <= 2230)) || ((pixel_index >= 2256) && (pixel_index <= 2257)) || ((pixel_index >= 2259) && (pixel_index <= 2264)) || ((pixel_index >= 2266) && (pixel_index <= 2267)) || ((pixel_index >= 2309) && (pixel_index <= 2326)) || ((pixel_index >= 2351) && (pixel_index <= 2360)) || ((pixel_index >= 2405) && (pixel_index <= 2422)) || ((pixel_index >= 2448) && (pixel_index <= 2459)) || ((pixel_index >= 2501) && (pixel_index <= 2518)) || ((pixel_index >= 2546) && (pixel_index <= 2556)) || ((pixel_index >= 2597) && (pixel_index <= 2614)) || ((pixel_index >= 2644) && (pixel_index <= 2652)) || ((pixel_index >= 2693) && (pixel_index <= 2710)) || ((pixel_index >= 2742) && (pixel_index <= 2750)) || ((pixel_index >= 2789) && (pixel_index <= 2806)) || ((pixel_index >= 2838) && (pixel_index <= 2846)) || ((pixel_index >= 2885) && (pixel_index <= 2902)) || ((pixel_index >= 2934) && (pixel_index <= 2938)) || ((pixel_index >= 2940) && (pixel_index <= 2941)) || ((pixel_index >= 2981) && (pixel_index <= 2998)) || ((pixel_index >= 3029) && (pixel_index <= 3034)) || ((pixel_index >= 3036) && (pixel_index <= 3037)) || ((pixel_index >= 3077) && (pixel_index <= 3094)) || ((pixel_index >= 3126) && (pixel_index <= 3133)) || ((pixel_index >= 3173) && (pixel_index <= 3190)) || ((pixel_index >= 3222) && (pixel_index <= 3230)) || ((pixel_index >= 3269) && (pixel_index <= 3286)) || ((pixel_index >= 3317) && (pixel_index <= 3318)) || ((pixel_index >= 3320) && (pixel_index <= 3328)) || ((pixel_index >= 3365) && (pixel_index <= 3382)) || ((pixel_index >= 3412) && (pixel_index <= 3413)) || ((pixel_index >= 3416) && (pixel_index <= 3427)) || ((pixel_index >= 3461) && (pixel_index <= 3478)) || ((pixel_index >= 3490) && (pixel_index <= 3494)) || pixel_index == 3508 || ((pixel_index >= 3510) && (pixel_index <= 3531)) || ((pixel_index >= 3557) && (pixel_index <= 3574)) || ((pixel_index >= 3587) && (pixel_index <= 3600)) || ((pixel_index >= 3602) && (pixel_index <= 3628)) || ((pixel_index >= 3653) && (pixel_index <= 3670)) || ((pixel_index >= 3686) && (pixel_index <= 3726)) || ((pixel_index >= 3749) && (pixel_index <= 3766)) || pixel_index == 3782 || ((pixel_index >= 3786) && (pixel_index <= 3788)) || ((pixel_index >= 3796) && (pixel_index <= 3822)) || ((pixel_index >= 3845) && (pixel_index <= 3862)) || ((pixel_index >= 3892) && (pixel_index <= 3919)) || ((pixel_index >= 3941) && (pixel_index <= 3958)) || ((pixel_index >= 3989) && (pixel_index <= 3997)) || ((pixel_index >= 4002) && (pixel_index <= 4014)) || ((pixel_index >= 4037) && (pixel_index <= 4054)) || ((pixel_index >= 4090) && (pixel_index <= 4093)) || ((pixel_index >= 4103) && (pixel_index <= 4108)) || ((pixel_index >= 4133) && (pixel_index <= 4150)) || ((pixel_index >= 4187) && (pixel_index <= 4189)) || ((pixel_index >= 4202) && (pixel_index <= 4203)) || ((pixel_index >= 4229) && (pixel_index <= 4246)) || ((pixel_index >= 4325) && (pixel_index <= 4342)) || ((pixel_index >= 4421) && (pixel_index <= 4438)) || ((pixel_index >= 4517) && (pixel_index <= 4534)) || ((pixel_index >= 4613) && (pixel_index <= 4630)) || ((pixel_index >= 4709) && (pixel_index <= 4726)) || ((pixel_index >= 4805) && (pixel_index <= 4822)) || ((pixel_index >= 4901) && (pixel_index <= 4918)) || ((pixel_index >= 4997) && (pixel_index <= 5014)) || ((pixel_index >= 5093) && (pixel_index <= 5110)) || ((pixel_index >= 5189) && (pixel_index <= 5206)) || ((pixel_index >= 5285) && (pixel_index <= 5302)) || ((pixel_index >= 5381) && (pixel_index <= 5398)) || ((pixel_index >= 5477) && (pixel_index <= 5494)) || ((pixel_index >= 5573) && (pixel_index <= 5590)) || ((pixel_index >= 5669) && (pixel_index <= 5686)) || ((pixel_index >= 5765) && (pixel_index <= 5782)) || ((pixel_index >= 5861) && (pixel_index <= 5878)) || ((pixel_index >= 5957) && (pixel_index <= 5974)) || (pixel_index >= 6053) && (pixel_index <= 6070)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 17) begin
            if (((pixel_index >= 5) && (pixel_index <= 19)) || ((pixel_index >= 101) && (pixel_index <= 115)) || ((pixel_index >= 197) && (pixel_index <= 211)) || ((pixel_index >= 293) && (pixel_index <= 307)) || ((pixel_index >= 389) && (pixel_index <= 403)) || ((pixel_index >= 485) && (pixel_index <= 499)) || ((pixel_index >= 581) && (pixel_index <= 595)) || ((pixel_index >= 677) && (pixel_index <= 691)) || ((pixel_index >= 773) && (pixel_index <= 787)) || ((pixel_index >= 869) && (pixel_index <= 883)) || ((pixel_index >= 965) && (pixel_index <= 979)) || ((pixel_index >= 1061) && (pixel_index <= 1075)) || ((pixel_index >= 1157) && (pixel_index <= 1171)) || ((pixel_index >= 1253) && (pixel_index <= 1267)) || ((pixel_index >= 1349) && (pixel_index <= 1363)) || ((pixel_index >= 1445) && (pixel_index <= 1459)) || ((pixel_index >= 1541) && (pixel_index <= 1555)) || ((pixel_index >= 1637) && (pixel_index <= 1651)) || ((pixel_index >= 1733) && (pixel_index <= 1747)) || ((pixel_index >= 1829) && (pixel_index <= 1843)) || ((pixel_index >= 1925) && (pixel_index <= 1939)) || ((pixel_index >= 2021) && (pixel_index <= 2035)) || ((pixel_index >= 2117) && (pixel_index <= 2131)) || ((pixel_index >= 2213) && (pixel_index <= 2227)) || pixel_index == 2262 || ((pixel_index >= 2309) && (pixel_index <= 2323)) || ((pixel_index >= 2352) && (pixel_index <= 2353)) || ((pixel_index >= 2356) && (pixel_index <= 2360)) || ((pixel_index >= 2405) && (pixel_index <= 2419)) || ((pixel_index >= 2447) && (pixel_index <= 2457)) || ((pixel_index >= 2501) && (pixel_index <= 2515)) || ((pixel_index >= 2543) && (pixel_index <= 2551)) || ((pixel_index >= 2553) && (pixel_index <= 2554)) || ((pixel_index >= 2597) && (pixel_index <= 2611)) || ((pixel_index >= 2641) && (pixel_index <= 2648)) || ((pixel_index >= 2693) && (pixel_index <= 2707)) || ((pixel_index >= 2738) && (pixel_index <= 2746)) || ((pixel_index >= 2789) && (pixel_index <= 2803)) || ((pixel_index >= 2836) && (pixel_index <= 2843)) || ((pixel_index >= 2885) && (pixel_index <= 2899)) || ((pixel_index >= 2933) && (pixel_index <= 2938)) || ((pixel_index >= 2981) && (pixel_index <= 2995)) || ((pixel_index >= 3029) && (pixel_index <= 3035)) || ((pixel_index >= 3077) && (pixel_index <= 3091)) || ((pixel_index >= 3124) && (pixel_index <= 3132)) || ((pixel_index >= 3173) && (pixel_index <= 3187)) || ((pixel_index >= 3220) && (pixel_index <= 3228)) || ((pixel_index >= 3269) && (pixel_index <= 3283)) || ((pixel_index >= 3317) && (pixel_index <= 3324)) || ((pixel_index >= 3365) && (pixel_index <= 3379)) || ((pixel_index >= 3413) && (pixel_index <= 3420)) || ((pixel_index >= 3461) && (pixel_index <= 3475)) || ((pixel_index >= 3508) && (pixel_index <= 3509)) || ((pixel_index >= 3511) && (pixel_index <= 3518)) || ((pixel_index >= 3557) && (pixel_index <= 3571)) || ((pixel_index >= 3586) && (pixel_index <= 3591)) || ((pixel_index >= 3603) && (pixel_index <= 3617)) || ((pixel_index >= 3621) && (pixel_index <= 3623)) || ((pixel_index >= 3653) && (pixel_index <= 3667)) || ((pixel_index >= 3683) && (pixel_index <= 3694)) || ((pixel_index >= 3698) && (pixel_index <= 3722)) || ((pixel_index >= 3749) && (pixel_index <= 3763)) || ((pixel_index >= 3781) && (pixel_index <= 3818)) || ((pixel_index >= 3845) && (pixel_index <= 3859)) || ((pixel_index >= 3881) && (pixel_index <= 3882)) || ((pixel_index >= 3890) && (pixel_index <= 3916)) || ((pixel_index >= 3941) && (pixel_index <= 3955)) || ((pixel_index >= 3978) && (pixel_index <= 3979)) || ((pixel_index >= 3987) && (pixel_index <= 4012)) || ((pixel_index >= 4037) && (pixel_index <= 4051)) || pixel_index == 4076 || ((pixel_index >= 4085) && (pixel_index <= 4108)) || ((pixel_index >= 4133) && (pixel_index <= 4147)) || ((pixel_index >= 4185) && (pixel_index <= 4188)) || ((pixel_index >= 4194) && (pixel_index <= 4204)) || ((pixel_index >= 4229) && (pixel_index <= 4243)) || ((pixel_index >= 4281) && (pixel_index <= 4284)) || ((pixel_index >= 4294) && (pixel_index <= 4298)) || ((pixel_index >= 4325) && (pixel_index <= 4339)) || ((pixel_index >= 4421) && (pixel_index <= 4435)) || ((pixel_index >= 4517) && (pixel_index <= 4531)) || ((pixel_index >= 4613) && (pixel_index <= 4627)) || ((pixel_index >= 4709) && (pixel_index <= 4723)) || ((pixel_index >= 4805) && (pixel_index <= 4819)) || ((pixel_index >= 4901) && (pixel_index <= 4915)) || ((pixel_index >= 4997) && (pixel_index <= 5011)) || ((pixel_index >= 5093) && (pixel_index <= 5107)) || ((pixel_index >= 5189) && (pixel_index <= 5203)) || ((pixel_index >= 5285) && (pixel_index <= 5299)) || ((pixel_index >= 5381) && (pixel_index <= 5395)) || ((pixel_index >= 5477) && (pixel_index <= 5491)) || ((pixel_index >= 5573) && (pixel_index <= 5587)) || ((pixel_index >= 5669) && (pixel_index <= 5683)) || ((pixel_index >= 5765) && (pixel_index <= 5779)) || ((pixel_index >= 5861) && (pixel_index <= 5875)) || ((pixel_index >= 5957) && (pixel_index <= 5971)) || (pixel_index >= 6053) && (pixel_index <= 6067)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 18) begin
            if (((pixel_index >= 5) && (pixel_index <= 21)) || ((pixel_index >= 101) && (pixel_index <= 117)) || ((pixel_index >= 197) && (pixel_index <= 213)) || ((pixel_index >= 293) && (pixel_index <= 309)) || ((pixel_index >= 389) && (pixel_index <= 405)) || ((pixel_index >= 485) && (pixel_index <= 501)) || ((pixel_index >= 581) && (pixel_index <= 597)) || ((pixel_index >= 677) && (pixel_index <= 693)) || ((pixel_index >= 773) && (pixel_index <= 789)) || ((pixel_index >= 869) && (pixel_index <= 885)) || ((pixel_index >= 965) && (pixel_index <= 981)) || ((pixel_index >= 1061) && (pixel_index <= 1077)) || ((pixel_index >= 1157) && (pixel_index <= 1173)) || ((pixel_index >= 1253) && (pixel_index <= 1269)) || ((pixel_index >= 1349) && (pixel_index <= 1365)) || ((pixel_index >= 1445) && (pixel_index <= 1461)) || ((pixel_index >= 1541) && (pixel_index <= 1557)) || ((pixel_index >= 1637) && (pixel_index <= 1653)) || ((pixel_index >= 1733) && (pixel_index <= 1749)) || ((pixel_index >= 1829) && (pixel_index <= 1845)) || ((pixel_index >= 1925) && (pixel_index <= 1941)) || ((pixel_index >= 2021) && (pixel_index <= 2037)) || ((pixel_index >= 2117) && (pixel_index <= 2133)) || ((pixel_index >= 2213) && (pixel_index <= 2229)) || ((pixel_index >= 2309) && (pixel_index <= 2325)) || ((pixel_index >= 2405) && (pixel_index <= 2421)) || ((pixel_index >= 2453) && (pixel_index <= 2455)) || ((pixel_index >= 2501) && (pixel_index <= 2517)) || ((pixel_index >= 2548) && (pixel_index <= 2551)) || ((pixel_index >= 2553) && (pixel_index <= 2557)) || ((pixel_index >= 2597) && (pixel_index <= 2613)) || ((pixel_index >= 2645) && (pixel_index <= 2654)) || ((pixel_index >= 2693) && (pixel_index <= 2709)) || ((pixel_index >= 2742) && (pixel_index <= 2751)) || ((pixel_index >= 2789) && (pixel_index <= 2805)) || ((pixel_index >= 2839) && (pixel_index <= 2844)) || pixel_index == 2847 || ((pixel_index >= 2885) && (pixel_index <= 2901)) || ((pixel_index >= 2935) && (pixel_index <= 2941)) || ((pixel_index >= 2981) && (pixel_index <= 2997)) || ((pixel_index >= 3032) && (pixel_index <= 3038)) || ((pixel_index >= 3077) && (pixel_index <= 3093)) || ((pixel_index >= 3129) && (pixel_index <= 3135)) || ((pixel_index >= 3173) && (pixel_index <= 3189)) || ((pixel_index >= 3225) && (pixel_index <= 3231)) || ((pixel_index >= 3269) && (pixel_index <= 3285)) || ((pixel_index >= 3321) && (pixel_index <= 3328)) || ((pixel_index >= 3365) && (pixel_index <= 3381)) || ((pixel_index >= 3416) && (pixel_index <= 3425)) || ((pixel_index >= 3461) && (pixel_index <= 3477)) || ((pixel_index >= 3513) && (pixel_index <= 3521)) || ((pixel_index >= 3557) && (pixel_index <= 3573)) || ((pixel_index >= 3609) && (pixel_index <= 3617)) || ((pixel_index >= 3653) && (pixel_index <= 3669)) || ((pixel_index >= 3686) && (pixel_index <= 3689)) || ((pixel_index >= 3704) && (pixel_index <= 3705)) || ((pixel_index >= 3707) && (pixel_index <= 3715)) || ((pixel_index >= 3749) && (pixel_index <= 3765)) || ((pixel_index >= 3783) && (pixel_index <= 3791)) || ((pixel_index >= 3799) && (pixel_index <= 3800)) || ((pixel_index >= 3802) && (pixel_index <= 3813)) || ((pixel_index >= 3845) && (pixel_index <= 3861)) || ((pixel_index >= 3881) && (pixel_index <= 3916)) || ((pixel_index >= 3941) && (pixel_index <= 3957)) || ((pixel_index >= 3981) && (pixel_index <= 4014)) || ((pixel_index >= 4037) && (pixel_index <= 4053)) || pixel_index == 4079 || ((pixel_index >= 4086) && (pixel_index <= 4111)) || ((pixel_index >= 4133) && (pixel_index <= 4149)) || ((pixel_index >= 4183) && (pixel_index <= 4208)) || ((pixel_index >= 4229) && (pixel_index <= 4245)) || ((pixel_index >= 4280) && (pixel_index <= 4305)) || ((pixel_index >= 4325) && (pixel_index <= 4341)) || ((pixel_index >= 4381) && (pixel_index <= 4383)) || ((pixel_index >= 4388) && (pixel_index <= 4401)) || ((pixel_index >= 4421) && (pixel_index <= 4437)) || ((pixel_index >= 4477) && (pixel_index <= 4479)) || ((pixel_index >= 4487) && (pixel_index <= 4496)) || ((pixel_index >= 4517) && (pixel_index <= 4533)) || pixel_index == 4573 || pixel_index == 4575 || ((pixel_index >= 4586) && (pixel_index <= 4590)) || pixel_index == 4592 || ((pixel_index >= 4613) && (pixel_index <= 4629)) || ((pixel_index >= 4684) && (pixel_index <= 4685)) || ((pixel_index >= 4709) && (pixel_index <= 4725)) || ((pixel_index >= 4805) && (pixel_index <= 4821)) || ((pixel_index >= 4901) && (pixel_index <= 4917)) || ((pixel_index >= 4997) && (pixel_index <= 5013)) || ((pixel_index >= 5093) && (pixel_index <= 5109)) || ((pixel_index >= 5189) && (pixel_index <= 5205)) || ((pixel_index >= 5285) && (pixel_index <= 5301)) || ((pixel_index >= 5381) && (pixel_index <= 5397)) || ((pixel_index >= 5477) && (pixel_index <= 5493)) || ((pixel_index >= 5573) && (pixel_index <= 5589)) || ((pixel_index >= 5669) && (pixel_index <= 5685)) || ((pixel_index >= 5765) && (pixel_index <= 5781)) || ((pixel_index >= 5861) && (pixel_index <= 5877)) || ((pixel_index >= 5957) && (pixel_index <= 5973)) || (pixel_index >= 6053) && (pixel_index <= 6069)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 19) begin
            if (((pixel_index >= 5) && (pixel_index <= 24)) || ((pixel_index >= 101) && (pixel_index <= 120)) || ((pixel_index >= 197) && (pixel_index <= 216)) || ((pixel_index >= 293) && (pixel_index <= 312)) || ((pixel_index >= 389) && (pixel_index <= 408)) || ((pixel_index >= 485) && (pixel_index <= 504)) || ((pixel_index >= 581) && (pixel_index <= 600)) || ((pixel_index >= 677) && (pixel_index <= 696)) || ((pixel_index >= 773) && (pixel_index <= 792)) || ((pixel_index >= 869) && (pixel_index <= 888)) || ((pixel_index >= 965) && (pixel_index <= 984)) || ((pixel_index >= 1061) && (pixel_index <= 1080)) || ((pixel_index >= 1157) && (pixel_index <= 1176)) || ((pixel_index >= 1253) && (pixel_index <= 1272)) || ((pixel_index >= 1349) && (pixel_index <= 1368)) || ((pixel_index >= 1445) && (pixel_index <= 1464)) || ((pixel_index >= 1541) && (pixel_index <= 1560)) || ((pixel_index >= 1637) && (pixel_index <= 1656)) || ((pixel_index >= 1733) && (pixel_index <= 1752)) || ((pixel_index >= 1829) && (pixel_index <= 1848)) || ((pixel_index >= 1925) && (pixel_index <= 1944)) || ((pixel_index >= 2021) && (pixel_index <= 2040)) || ((pixel_index >= 2117) && (pixel_index <= 2136)) || ((pixel_index >= 2213) && (pixel_index <= 2232)) || pixel_index == 2267 || ((pixel_index >= 2309) && (pixel_index <= 2328)) || ((pixel_index >= 2362) && (pixel_index <= 2364)) || ((pixel_index >= 2405) && (pixel_index <= 2424)) || ((pixel_index >= 2458) && (pixel_index <= 2460)) || pixel_index == 2464 || ((pixel_index >= 2501) && (pixel_index <= 2520)) || ((pixel_index >= 2554) && (pixel_index <= 2562)) || ((pixel_index >= 2597) && (pixel_index <= 2616)) || ((pixel_index >= 2651) && (pixel_index <= 2659)) || ((pixel_index >= 2693) && (pixel_index <= 2712)) || ((pixel_index >= 2748) && (pixel_index <= 2756)) || ((pixel_index >= 2790) && (pixel_index <= 2808)) || ((pixel_index >= 2844) && (pixel_index <= 2849)) || ((pixel_index >= 2852) && (pixel_index <= 2853)) || ((pixel_index >= 2886) && (pixel_index <= 2904)) || ((pixel_index >= 2940) && (pixel_index <= 2945)) || pixel_index == 2949 || ((pixel_index >= 2982) && (pixel_index <= 3000)) || ((pixel_index >= 3037) && (pixel_index <= 3042)) || ((pixel_index >= 3078) && (pixel_index <= 3096)) || ((pixel_index >= 3133) && (pixel_index <= 3139)) || ((pixel_index >= 3174) && (pixel_index <= 3192)) || ((pixel_index >= 3229) && (pixel_index <= 3235)) || ((pixel_index >= 3269) && (pixel_index <= 3288)) || ((pixel_index >= 3324) && (pixel_index <= 3332)) || ((pixel_index >= 3365) && (pixel_index <= 3384)) || ((pixel_index >= 3421) && (pixel_index <= 3429)) || ((pixel_index >= 3461) && (pixel_index <= 3480)) || ((pixel_index >= 3497) && (pixel_index <= 3499)) || ((pixel_index >= 3517) && (pixel_index <= 3525)) || ((pixel_index >= 3557) && (pixel_index <= 3576)) || ((pixel_index >= 3594) && (pixel_index <= 3598)) || ((pixel_index >= 3612) && (pixel_index <= 3613)) || ((pixel_index >= 3615) && (pixel_index <= 3620)) || ((pixel_index >= 3653) && (pixel_index <= 3672)) || ((pixel_index >= 3692) && (pixel_index <= 3698)) || ((pixel_index >= 3707) && (pixel_index <= 3709)) || ((pixel_index >= 3711) && (pixel_index <= 3717)) || ((pixel_index >= 3749) && (pixel_index <= 3768)) || ((pixel_index >= 3788) && (pixel_index <= 3797)) || ((pixel_index >= 3802) && (pixel_index <= 3804)) || ((pixel_index >= 3806) && (pixel_index <= 3814)) || ((pixel_index >= 3845) && (pixel_index <= 3864)) || pixel_index == 3888 || ((pixel_index >= 3891) && (pixel_index <= 3908)) || ((pixel_index >= 3910) && (pixel_index <= 3914)) || ((pixel_index >= 3941) && (pixel_index <= 3960)) || pixel_index == 3985 || ((pixel_index >= 3991) && (pixel_index <= 4005)) || ((pixel_index >= 4008) && (pixel_index <= 4009)) || ((pixel_index >= 4037) && (pixel_index <= 4056)) || ((pixel_index >= 4082) && (pixel_index <= 4083)) || ((pixel_index >= 4090) && (pixel_index <= 4112)) || ((pixel_index >= 4133) && (pixel_index <= 4152)) || ((pixel_index >= 4186) && (pixel_index <= 4210)) || ((pixel_index >= 4229) && (pixel_index <= 4248)) || ((pixel_index >= 4283) && (pixel_index <= 4307)) || ((pixel_index >= 4325) && (pixel_index <= 4344)) || ((pixel_index >= 4383) && (pixel_index <= 4404)) || ((pixel_index >= 4421) && (pixel_index <= 4440)) || ((pixel_index >= 4480) && (pixel_index <= 4501)) || ((pixel_index >= 4517) && (pixel_index <= 4536)) || ((pixel_index >= 4576) && (pixel_index <= 4579)) || ((pixel_index >= 4584) && (pixel_index <= 4597)) || ((pixel_index >= 4613) && (pixel_index <= 4632)) || ((pixel_index >= 4672) && (pixel_index <= 4675)) || ((pixel_index >= 4683) && (pixel_index <= 4693)) || ((pixel_index >= 4709) && (pixel_index <= 4728)) || ((pixel_index >= 4781) && (pixel_index <= 4788)) || ((pixel_index >= 4805) && (pixel_index <= 4824)) || ((pixel_index >= 4879) && (pixel_index <= 4882)) || ((pixel_index >= 4901) && (pixel_index <= 4920)) || ((pixel_index >= 4997) && (pixel_index <= 5016)) || ((pixel_index >= 5093) && (pixel_index <= 5112)) || ((pixel_index >= 5189) && (pixel_index <= 5208)) || ((pixel_index >= 5285) && (pixel_index <= 5304)) || ((pixel_index >= 5381) && (pixel_index <= 5400)) || ((pixel_index >= 5477) && (pixel_index <= 5496)) || ((pixel_index >= 5573) && (pixel_index <= 5592)) || ((pixel_index >= 5669) && (pixel_index <= 5688)) || ((pixel_index >= 5765) && (pixel_index <= 5784)) || ((pixel_index >= 5861) && (pixel_index <= 5880)) || ((pixel_index >= 5957) && (pixel_index <= 5976)) || (pixel_index >= 6053) && (pixel_index <= 6072)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 20) begin
            if (((pixel_index >= 5) && (pixel_index <= 28)) || ((pixel_index >= 101) && (pixel_index <= 124)) || ((pixel_index >= 197) && (pixel_index <= 220)) || ((pixel_index >= 293) && (pixel_index <= 316)) || ((pixel_index >= 389) && (pixel_index <= 412)) || ((pixel_index >= 485) && (pixel_index <= 508)) || ((pixel_index >= 581) && (pixel_index <= 604)) || ((pixel_index >= 677) && (pixel_index <= 700)) || ((pixel_index >= 773) && (pixel_index <= 796)) || ((pixel_index >= 869) && (pixel_index <= 892)) || ((pixel_index >= 965) && (pixel_index <= 988)) || ((pixel_index >= 1061) && (pixel_index <= 1084)) || ((pixel_index >= 1157) && (pixel_index <= 1180)) || ((pixel_index >= 1253) && (pixel_index <= 1276)) || ((pixel_index >= 1349) && (pixel_index <= 1372)) || ((pixel_index >= 1445) && (pixel_index <= 1468)) || ((pixel_index >= 1541) && (pixel_index <= 1564)) || ((pixel_index >= 1637) && (pixel_index <= 1660)) || ((pixel_index >= 1733) && (pixel_index <= 1756)) || ((pixel_index >= 1791) && (pixel_index <= 1792)) || ((pixel_index >= 1829) && (pixel_index <= 1852)) || ((pixel_index >= 1886) && (pixel_index <= 1888)) || ((pixel_index >= 1925) && (pixel_index <= 1948)) || ((pixel_index >= 1982) && (pixel_index <= 1984)) || pixel_index == 1988 || ((pixel_index >= 2021) && (pixel_index <= 2044)) || ((pixel_index >= 2079) && (pixel_index <= 2086)) || ((pixel_index >= 2117) && (pixel_index <= 2140)) || ((pixel_index >= 2175) && (pixel_index <= 2182)) || ((pixel_index >= 2213) && (pixel_index <= 2236)) || ((pixel_index >= 2272) && (pixel_index <= 2279)) || ((pixel_index >= 2309) && (pixel_index <= 2332)) || ((pixel_index >= 2368) && (pixel_index <= 2375)) || ((pixel_index >= 2407) && (pixel_index <= 2428)) || ((pixel_index >= 2464) && (pixel_index <= 2469)) || ((pixel_index >= 2471) && (pixel_index <= 2472)) || ((pixel_index >= 2504) && (pixel_index <= 2524)) || ((pixel_index >= 2561) && (pixel_index <= 2565)) || pixel_index == 2568 || ((pixel_index >= 2601) && (pixel_index <= 2620)) || ((pixel_index >= 2657) && (pixel_index <= 2661)) || ((pixel_index >= 2697) && (pixel_index <= 2716)) || ((pixel_index >= 2752) && (pixel_index <= 2756)) || pixel_index == 2758 || ((pixel_index >= 2794) && (pixel_index <= 2812)) || pixel_index == 2828 || ((pixel_index >= 2848) && (pixel_index <= 2854)) || ((pixel_index >= 2890) && (pixel_index <= 2908)) || ((pixel_index >= 2924) && (pixel_index <= 2927)) || ((pixel_index >= 2944) && (pixel_index <= 2949)) || ((pixel_index >= 2986) && (pixel_index <= 3004)) || ((pixel_index >= 3020) && (pixel_index <= 3025)) || ((pixel_index >= 3039) && (pixel_index <= 3045)) || ((pixel_index >= 3082) && (pixel_index <= 3100)) || ((pixel_index >= 3118) && (pixel_index <= 3124)) || ((pixel_index >= 3135) && (pixel_index <= 3136)) || ((pixel_index >= 3138) && (pixel_index <= 3143)) || ((pixel_index >= 3178) && (pixel_index <= 3196)) || ((pixel_index >= 3214) && (pixel_index <= 3222)) || ((pixel_index >= 3230) && (pixel_index <= 3232)) || ((pixel_index >= 3234) && (pixel_index <= 3239)) || ((pixel_index >= 3273) && (pixel_index <= 3292)) || ((pixel_index >= 3314) && (pixel_index <= 3321)) || ((pixel_index >= 3324) && (pixel_index <= 3326)) || ((pixel_index >= 3329) && (pixel_index <= 3335)) || ((pixel_index >= 3369) && (pixel_index <= 3388)) || pixel_index == 3411 || ((pixel_index >= 3415) && (pixel_index <= 3432)) || ((pixel_index >= 3464) && (pixel_index <= 3484)) || ((pixel_index >= 3507) && (pixel_index <= 3508)) || ((pixel_index >= 3514) && (pixel_index <= 3529)) || ((pixel_index >= 3559) && (pixel_index <= 3580)) || ((pixel_index >= 3603) && (pixel_index <= 3604)) || ((pixel_index >= 3612) && (pixel_index <= 3626)) || ((pixel_index >= 3653) && (pixel_index <= 3676)) || pixel_index == 3700 || ((pixel_index >= 3709) && (pixel_index <= 3727)) || ((pixel_index >= 3749) && (pixel_index <= 3772)) || ((pixel_index >= 3805) && (pixel_index <= 3827)) || ((pixel_index >= 3845) && (pixel_index <= 3868)) || ((pixel_index >= 3903) && (pixel_index <= 3925)) || ((pixel_index >= 3941) && (pixel_index <= 3964)) || ((pixel_index >= 4001) && (pixel_index <= 4021)) || ((pixel_index >= 4037) && (pixel_index <= 4060)) || ((pixel_index >= 4098) && (pixel_index <= 4118)) || ((pixel_index >= 4133) && (pixel_index <= 4156)) || ((pixel_index >= 4194) && (pixel_index <= 4198)) || ((pixel_index >= 4202) && (pixel_index <= 4215)) || ((pixel_index >= 4229) && (pixel_index <= 4252)) || ((pixel_index >= 4291) && (pixel_index <= 4293)) || ((pixel_index >= 4300) && (pixel_index <= 4311)) || ((pixel_index >= 4325) && (pixel_index <= 4348)) || ((pixel_index >= 4398) && (pixel_index <= 4407)) || ((pixel_index >= 4421) && (pixel_index <= 4444)) || ((pixel_index >= 4496) && (pixel_index <= 4503)) || ((pixel_index >= 4517) && (pixel_index <= 4540)) || ((pixel_index >= 4593) && (pixel_index <= 4599)) || ((pixel_index >= 4613) && (pixel_index <= 4636)) || pixel_index == 4691 || ((pixel_index >= 4709) && (pixel_index <= 4732)) || ((pixel_index >= 4805) && (pixel_index <= 4828)) || ((pixel_index >= 4901) && (pixel_index <= 4924)) || ((pixel_index >= 4997) && (pixel_index <= 5020)) || ((pixel_index >= 5093) && (pixel_index <= 5116)) || ((pixel_index >= 5189) && (pixel_index <= 5212)) || ((pixel_index >= 5285) && (pixel_index <= 5308)) || ((pixel_index >= 5381) && (pixel_index <= 5404)) || ((pixel_index >= 5477) && (pixel_index <= 5500)) || ((pixel_index >= 5573) && (pixel_index <= 5596)) || ((pixel_index >= 5669) && (pixel_index <= 5692)) || ((pixel_index >= 5765) && (pixel_index <= 5788)) || ((pixel_index >= 5861) && (pixel_index <= 5884)) || ((pixel_index >= 5957) && (pixel_index <= 5980)) || (pixel_index >= 6053) && (pixel_index <= 6076)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 21) begin
            if (((pixel_index >= 5) && (pixel_index <= 40)) || ((pixel_index >= 70) && (pixel_index <= 79)) || ((pixel_index >= 101) && (pixel_index <= 137)) || ((pixel_index >= 167) && (pixel_index <= 176)) || ((pixel_index >= 197) && (pixel_index <= 233)) || ((pixel_index >= 263) && (pixel_index <= 272)) || ((pixel_index >= 293) && (pixel_index <= 328)) || ((pixel_index >= 360) && (pixel_index <= 368)) || ((pixel_index >= 389) && (pixel_index <= 425)) || ((pixel_index >= 457) && (pixel_index <= 464)) || ((pixel_index >= 485) && (pixel_index <= 520)) || ((pixel_index >= 553) && (pixel_index <= 561)) || ((pixel_index >= 581) && (pixel_index <= 616)) || ((pixel_index >= 650) && (pixel_index <= 656)) || ((pixel_index >= 677) && (pixel_index <= 712)) || ((pixel_index >= 746) && (pixel_index <= 752)) || ((pixel_index >= 773) && (pixel_index <= 808)) || ((pixel_index >= 841) && (pixel_index <= 849)) || ((pixel_index >= 869) && (pixel_index <= 904)) || ((pixel_index >= 937) && (pixel_index <= 944)) || ((pixel_index >= 965) && (pixel_index <= 1000)) || ((pixel_index >= 1012) && (pixel_index <= 1014)) || ((pixel_index >= 1033) && (pixel_index <= 1040)) || ((pixel_index >= 1061) && (pixel_index <= 1096)) || ((pixel_index >= 1109) && (pixel_index <= 1112)) || ((pixel_index >= 1128) && (pixel_index <= 1136)) || ((pixel_index >= 1157) && (pixel_index <= 1192)) || ((pixel_index >= 1205) && (pixel_index <= 1211)) || ((pixel_index >= 1224) && (pixel_index <= 1232)) || ((pixel_index >= 1253) && (pixel_index <= 1288)) || ((pixel_index >= 1303) && (pixel_index <= 1310)) || ((pixel_index >= 1319) && (pixel_index <= 1328)) || ((pixel_index >= 1349) && (pixel_index <= 1384)) || ((pixel_index >= 1400) && (pixel_index <= 1409)) || ((pixel_index >= 1414) && (pixel_index <= 1425)) || ((pixel_index >= 1445) && (pixel_index <= 1480)) || ((pixel_index >= 1499) && (pixel_index <= 1522)) || ((pixel_index >= 1541) && (pixel_index <= 1576)) || ((pixel_index >= 1596) && (pixel_index <= 1619)) || ((pixel_index >= 1637) && (pixel_index <= 1672)) || ((pixel_index >= 1694) && (pixel_index <= 1695)) || ((pixel_index >= 1698) && (pixel_index <= 1716)) || ((pixel_index >= 1733) && (pixel_index <= 1768)) || ((pixel_index >= 1797) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1864)) || ((pixel_index >= 1894) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 1960)) || ((pixel_index >= 1990) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2056)) || ((pixel_index >= 2089) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2152)) || ((pixel_index >= 2187) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2248)) || ((pixel_index >= 2284) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2316)) || ((pixel_index >= 2321) && (pixel_index <= 2344)) || ((pixel_index >= 2380) && (pixel_index <= 2382)) || ((pixel_index >= 2388) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2410)) || ((pixel_index >= 2419) && (pixel_index <= 2440)) || ((pixel_index >= 2476) && (pixel_index <= 2477)) || ((pixel_index >= 2486) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2505)) || ((pixel_index >= 2516) && (pixel_index <= 2536)) || ((pixel_index >= 2584) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2600)) || ((pixel_index >= 2613) && (pixel_index <= 2632)) || ((pixel_index >= 2693) && (pixel_index <= 2696)) || ((pixel_index >= 2709) && (pixel_index <= 2728)) || ((pixel_index >= 2789) && (pixel_index <= 2791)) || ((pixel_index >= 2806) && (pixel_index <= 2824)) || ((pixel_index >= 2885) && (pixel_index <= 2887)) || ((pixel_index >= 2902) && (pixel_index <= 2920)) || ((pixel_index >= 2981) && (pixel_index <= 2983)) || ((pixel_index >= 2998) && (pixel_index <= 3016)) || ((pixel_index >= 3077) && (pixel_index <= 3079)) || ((pixel_index >= 3094) && (pixel_index <= 3112)) || ((pixel_index >= 3173) && (pixel_index <= 3175)) || ((pixel_index >= 3190) && (pixel_index <= 3208)) || ((pixel_index >= 3269) && (pixel_index <= 3272)) || ((pixel_index >= 3285) && (pixel_index <= 3304)) || ((pixel_index >= 3365) && (pixel_index <= 3368)) || ((pixel_index >= 3381) && (pixel_index <= 3400)) || ((pixel_index >= 3461) && (pixel_index <= 3465)) || ((pixel_index >= 3476) && (pixel_index <= 3496)) || ((pixel_index >= 3557) && (pixel_index <= 3562)) || ((pixel_index >= 3571) && (pixel_index <= 3592)) || ((pixel_index >= 3653) && (pixel_index <= 3660)) || ((pixel_index >= 3665) && (pixel_index <= 3688)) || ((pixel_index >= 3749) && (pixel_index <= 3784)) || ((pixel_index >= 3845) && (pixel_index <= 3880)) || ((pixel_index >= 3941) && (pixel_index <= 3976)) || ((pixel_index >= 4037) && (pixel_index <= 4072)) || ((pixel_index >= 4133) && (pixel_index <= 4168)) || ((pixel_index >= 4229) && (pixel_index <= 4264)) || ((pixel_index >= 4325) && (pixel_index <= 4360)) || ((pixel_index >= 4421) && (pixel_index <= 4456)) || ((pixel_index >= 4517) && (pixel_index <= 4552)) || ((pixel_index >= 4613) && (pixel_index <= 4648)) || ((pixel_index >= 4709) && (pixel_index <= 4744)) || ((pixel_index >= 4805) && (pixel_index <= 4840)) || ((pixel_index >= 4901) && (pixel_index <= 4936)) || ((pixel_index >= 4997) && (pixel_index <= 5032)) || ((pixel_index >= 5093) && (pixel_index <= 5128)) || ((pixel_index >= 5189) && (pixel_index <= 5224)) || ((pixel_index >= 5285) && (pixel_index <= 5320)) || ((pixel_index >= 5381) && (pixel_index <= 5416)) || ((pixel_index >= 5477) && (pixel_index <= 5512)) || ((pixel_index >= 5573) && (pixel_index <= 5608)) || ((pixel_index >= 5669) && (pixel_index <= 5704)) || ((pixel_index >= 5765) && (pixel_index <= 5800)) || ((pixel_index >= 5861) && (pixel_index <= 5896)) || ((pixel_index >= 5957) && (pixel_index <= 5992)) || (pixel_index >= 6053) && (pixel_index <= 6088)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 22) begin
            if (((pixel_index >= 5) && (pixel_index <= 68)) || ((pixel_index >= 101) && (pixel_index <= 164)) || ((pixel_index >= 197) && (pixel_index <= 260)) || ((pixel_index >= 293) && (pixel_index <= 356)) || ((pixel_index >= 389) && (pixel_index <= 452)) || ((pixel_index >= 485) && (pixel_index <= 548)) || ((pixel_index >= 581) && (pixel_index <= 644)) || ((pixel_index >= 677) && (pixel_index <= 740)) || ((pixel_index >= 773) && (pixel_index <= 836)) || ((pixel_index >= 869) && (pixel_index <= 932)) || ((pixel_index >= 965) && (pixel_index <= 1028)) || ((pixel_index >= 1061) && (pixel_index <= 1124)) || ((pixel_index >= 1157) && (pixel_index <= 1220)) || ((pixel_index >= 1253) && (pixel_index <= 1316)) || ((pixel_index >= 1349) && (pixel_index <= 1412)) || ((pixel_index >= 1445) && (pixel_index <= 1508)) || ((pixel_index >= 1541) && (pixel_index <= 1604)) || ((pixel_index >= 1637) && (pixel_index <= 1700)) || ((pixel_index >= 1733) && (pixel_index <= 1796)) || ((pixel_index >= 1829) && (pixel_index <= 1892)) || ((pixel_index >= 1925) && (pixel_index <= 1988)) || ((pixel_index >= 2021) && (pixel_index <= 2053)) || pixel_index == 2055 || ((pixel_index >= 2057) && (pixel_index <= 2084)) || ((pixel_index >= 2117) && (pixel_index <= 2147)) || ((pixel_index >= 2157) && (pixel_index <= 2180)) || ((pixel_index >= 2213) && (pixel_index <= 2241)) || ((pixel_index >= 2254) && (pixel_index <= 2276)) || ((pixel_index >= 2309) && (pixel_index <= 2336)) || ((pixel_index >= 2351) && (pixel_index <= 2372)) || ((pixel_index >= 2405) && (pixel_index <= 2431)) || ((pixel_index >= 2447) && (pixel_index <= 2468)) || ((pixel_index >= 2501) && (pixel_index <= 2526)) || ((pixel_index >= 2544) && (pixel_index <= 2564)) || ((pixel_index >= 2597) && (pixel_index <= 2622)) || ((pixel_index >= 2640) && (pixel_index <= 2660)) || ((pixel_index >= 2693) && (pixel_index <= 2718)) || ((pixel_index >= 2736) && (pixel_index <= 2756)) || ((pixel_index >= 2789) && (pixel_index <= 2814)) || ((pixel_index >= 2832) && (pixel_index <= 2852)) || ((pixel_index >= 2885) && (pixel_index <= 2910)) || ((pixel_index >= 2928) && (pixel_index <= 2948)) || ((pixel_index >= 2981) && (pixel_index <= 3007)) || ((pixel_index >= 3024) && (pixel_index <= 3044)) || ((pixel_index >= 3077) && (pixel_index <= 3103)) || ((pixel_index >= 3120) && (pixel_index <= 3140)) || ((pixel_index >= 3173) && (pixel_index <= 3199)) || ((pixel_index >= 3215) && (pixel_index <= 3236)) || ((pixel_index >= 3269) && (pixel_index <= 3296)) || ((pixel_index >= 3311) && (pixel_index <= 3332)) || ((pixel_index >= 3365) && (pixel_index <= 3393)) || ((pixel_index >= 3406) && (pixel_index <= 3428)) || ((pixel_index >= 3461) && (pixel_index <= 3489)) || ((pixel_index >= 3501) && (pixel_index <= 3524)) || ((pixel_index >= 3557) && (pixel_index <= 3587)) || ((pixel_index >= 3596) && (pixel_index <= 3620)) || ((pixel_index >= 3653) && (pixel_index <= 3685)) || ((pixel_index >= 3690) && (pixel_index <= 3716)) || ((pixel_index >= 3749) && (pixel_index <= 3812)) || ((pixel_index >= 3845) && (pixel_index <= 3908)) || ((pixel_index >= 3941) && (pixel_index <= 4004)) || ((pixel_index >= 4037) && (pixel_index <= 4100)) || ((pixel_index >= 4133) && (pixel_index <= 4196)) || ((pixel_index >= 4229) && (pixel_index <= 4292)) || ((pixel_index >= 4325) && (pixel_index <= 4388)) || ((pixel_index >= 4421) && (pixel_index <= 4484)) || ((pixel_index >= 4517) && (pixel_index <= 4580)) || ((pixel_index >= 4613) && (pixel_index <= 4676)) || ((pixel_index >= 4709) && (pixel_index <= 4772)) || ((pixel_index >= 4805) && (pixel_index <= 4868)) || ((pixel_index >= 4901) && (pixel_index <= 4964)) || ((pixel_index >= 4997) && (pixel_index <= 5060)) || ((pixel_index >= 5093) && (pixel_index <= 5156)) || ((pixel_index >= 5189) && (pixel_index <= 5252)) || ((pixel_index >= 5285) && (pixel_index <= 5348)) || ((pixel_index >= 5381) && (pixel_index <= 5444)) || ((pixel_index >= 5477) && (pixel_index <= 5540)) || ((pixel_index >= 5573) && (pixel_index <= 5636)) || ((pixel_index >= 5669) && (pixel_index <= 5732)) || ((pixel_index >= 5765) && (pixel_index <= 5828)) || ((pixel_index >= 5861) && (pixel_index <= 5924)) || ((pixel_index >= 5957) && (pixel_index <= 6020)) || (pixel_index >= 6053) && (pixel_index <= 6116)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 23) begin
            if (((pixel_index >= 5) && (pixel_index <= 87)) || ((pixel_index >= 101) && (pixel_index <= 183)) || ((pixel_index >= 197) && (pixel_index <= 279)) || ((pixel_index >= 293) && (pixel_index <= 375)) || ((pixel_index >= 389) && (pixel_index <= 471)) || ((pixel_index >= 485) && (pixel_index <= 567)) || ((pixel_index >= 581) && (pixel_index <= 663)) || ((pixel_index >= 677) && (pixel_index <= 759)) || ((pixel_index >= 773) && (pixel_index <= 855)) || ((pixel_index >= 869) && (pixel_index <= 951)) || ((pixel_index >= 965) && (pixel_index <= 1047)) || ((pixel_index >= 1061) && (pixel_index <= 1143)) || ((pixel_index >= 1157) && (pixel_index <= 1239)) || ((pixel_index >= 1253) && (pixel_index <= 1335)) || ((pixel_index >= 1349) && (pixel_index <= 1431)) || ((pixel_index >= 1445) && (pixel_index <= 1527)) || ((pixel_index >= 1541) && (pixel_index <= 1623)) || ((pixel_index >= 1637) && (pixel_index <= 1680)) || ((pixel_index >= 1682) && (pixel_index <= 1719)) || ((pixel_index >= 1733) && (pixel_index <= 1776)) || ((pixel_index >= 1778) && (pixel_index <= 1815)) || ((pixel_index >= 1829) && (pixel_index <= 1867)) || ((pixel_index >= 1874) && (pixel_index <= 1911)) || ((pixel_index >= 1925) && (pixel_index <= 1961)) || ((pixel_index >= 1974) && (pixel_index <= 2007)) || ((pixel_index >= 2021) && (pixel_index <= 2056)) || ((pixel_index >= 2072) && (pixel_index <= 2103)) || ((pixel_index >= 2117) && (pixel_index <= 2151)) || ((pixel_index >= 2168) && (pixel_index <= 2199)) || ((pixel_index >= 2213) && (pixel_index <= 2247)) || ((pixel_index >= 2265) && (pixel_index <= 2295)) || ((pixel_index >= 2309) && (pixel_index <= 2343)) || ((pixel_index >= 2361) && (pixel_index <= 2391)) || ((pixel_index >= 2405) && (pixel_index <= 2439)) || ((pixel_index >= 2458) && (pixel_index <= 2487)) || ((pixel_index >= 2501) && (pixel_index <= 2534)) || ((pixel_index >= 2554) && (pixel_index <= 2583)) || ((pixel_index >= 2597) && (pixel_index <= 2630)) || ((pixel_index >= 2650) && (pixel_index <= 2679)) || ((pixel_index >= 2693) && (pixel_index <= 2727)) || ((pixel_index >= 2745) && (pixel_index <= 2775)) || ((pixel_index >= 2789) && (pixel_index <= 2823)) || ((pixel_index >= 2841) && (pixel_index <= 2871)) || ((pixel_index >= 2885) && (pixel_index <= 2919)) || ((pixel_index >= 2937) && (pixel_index <= 2967)) || ((pixel_index >= 2981) && (pixel_index <= 3015)) || ((pixel_index >= 3033) && (pixel_index <= 3063)) || ((pixel_index >= 3077) && (pixel_index <= 3112)) || ((pixel_index >= 3128) && (pixel_index <= 3159)) || ((pixel_index >= 3173) && (pixel_index <= 3208)) || ((pixel_index >= 3223) && (pixel_index <= 3255)) || ((pixel_index >= 3269) && (pixel_index <= 3305)) || ((pixel_index >= 3319) && (pixel_index <= 3351)) || ((pixel_index >= 3365) && (pixel_index <= 3402)) || ((pixel_index >= 3414) && (pixel_index <= 3447)) || ((pixel_index >= 3461) && (pixel_index <= 3499)) || pixel_index == 3503 || ((pixel_index >= 3508) && (pixel_index <= 3543)) || ((pixel_index >= 3557) && (pixel_index <= 3639)) || ((pixel_index >= 3653) && (pixel_index <= 3735)) || ((pixel_index >= 3749) && (pixel_index <= 3831)) || ((pixel_index >= 3845) && (pixel_index <= 3927)) || ((pixel_index >= 3941) && (pixel_index <= 4023)) || ((pixel_index >= 4037) && (pixel_index <= 4119)) || ((pixel_index >= 4133) && (pixel_index <= 4215)) || ((pixel_index >= 4229) && (pixel_index <= 4311)) || ((pixel_index >= 4325) && (pixel_index <= 4407)) || ((pixel_index >= 4421) && (pixel_index <= 4503)) || ((pixel_index >= 4517) && (pixel_index <= 4599)) || ((pixel_index >= 4613) && (pixel_index <= 4695)) || ((pixel_index >= 4709) && (pixel_index <= 4791)) || ((pixel_index >= 4805) && (pixel_index <= 4887)) || ((pixel_index >= 4901) && (pixel_index <= 4983)) || ((pixel_index >= 4997) && (pixel_index <= 5079)) || ((pixel_index >= 5093) && (pixel_index <= 5175)) || ((pixel_index >= 5189) && (pixel_index <= 5271)) || ((pixel_index >= 5285) && (pixel_index <= 5367)) || ((pixel_index >= 5381) && (pixel_index <= 5463)) || ((pixel_index >= 5477) && (pixel_index <= 5559)) || ((pixel_index >= 5573) && (pixel_index <= 5655)) || ((pixel_index >= 5669) && (pixel_index <= 5751)) || ((pixel_index >= 5765) && (pixel_index <= 5847)) || ((pixel_index >= 5861) && (pixel_index <= 5943)) || ((pixel_index >= 5957) && (pixel_index <= 6039)) || (pixel_index >= 6053) && (pixel_index <= 6135)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 24) begin
            if (((pixel_index >= 8) && (pixel_index <= 89)) || ((pixel_index >= 103) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 377)) || ((pixel_index >= 389) && (pixel_index <= 473)) || ((pixel_index >= 485) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 857)) || ((pixel_index >= 869) && (pixel_index <= 953)) || ((pixel_index >= 965) && (pixel_index <= 1049)) || ((pixel_index >= 1061) && (pixel_index <= 1145)) || ((pixel_index >= 1157) && (pixel_index <= 1241)) || ((pixel_index >= 1254) && (pixel_index <= 1337)) || ((pixel_index >= 1350) && (pixel_index <= 1433)) || ((pixel_index >= 1446) && (pixel_index <= 1529)) || ((pixel_index >= 1541) && (pixel_index <= 1625)) || ((pixel_index >= 1637) && (pixel_index <= 1721)) || ((pixel_index >= 1733) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2639)) || ((pixel_index >= 2647) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2734)) || ((pixel_index >= 2745) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2830)) || ((pixel_index >= 2843) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2925)) || ((pixel_index >= 2939) && (pixel_index <= 2969)) || ((pixel_index >= 2982) && (pixel_index <= 3021)) || ((pixel_index >= 3036) && (pixel_index <= 3065)) || ((pixel_index >= 3079) && (pixel_index <= 3116)) || ((pixel_index >= 3133) && (pixel_index <= 3161)) || ((pixel_index >= 3175) && (pixel_index <= 3212)) || ((pixel_index >= 3229) && (pixel_index <= 3257)) || ((pixel_index >= 3271) && (pixel_index <= 3308)) || ((pixel_index >= 3326) && (pixel_index <= 3353)) || ((pixel_index >= 3368) && (pixel_index <= 3404)) || ((pixel_index >= 3422) && (pixel_index <= 3449)) || ((pixel_index >= 3464) && (pixel_index <= 3500)) || ((pixel_index >= 3518) && (pixel_index <= 3545)) || ((pixel_index >= 3562) && (pixel_index <= 3581)) || ((pixel_index >= 3592) && (pixel_index <= 3596)) || ((pixel_index >= 3614) && (pixel_index <= 3641)) || ((pixel_index >= 3659) && (pixel_index <= 3662)) || ((pixel_index >= 3689) && (pixel_index <= 3691)) || ((pixel_index >= 3710) && (pixel_index <= 3737)) || ((pixel_index >= 3805) && (pixel_index <= 3833)) || ((pixel_index >= 3901) && (pixel_index <= 3929)) || ((pixel_index >= 3997) && (pixel_index <= 4025)) || ((pixel_index >= 4092) && (pixel_index <= 4121)) || ((pixel_index >= 4188) && (pixel_index <= 4217)) || ((pixel_index >= 4282) && (pixel_index <= 4313)) || ((pixel_index >= 4377) && (pixel_index <= 4409)) || pixel_index == 4460 || ((pixel_index >= 4472) && (pixel_index <= 4505)) || ((pixel_index >= 4555) && (pixel_index <= 4560)) || ((pixel_index >= 4563) && (pixel_index <= 4564)) || ((pixel_index >= 4566) && (pixel_index <= 4601)) || ((pixel_index >= 4651) && (pixel_index <= 4697)) || ((pixel_index >= 4748) && (pixel_index <= 4793)) || ((pixel_index >= 4844) && (pixel_index <= 4889)) || ((pixel_index >= 4940) && (pixel_index <= 4985)) || ((pixel_index >= 5036) && (pixel_index <= 5081)) || ((pixel_index >= 5132) && (pixel_index <= 5177)) || ((pixel_index >= 5228) && (pixel_index <= 5273)) || ((pixel_index >= 5325) && (pixel_index <= 5369)) || ((pixel_index >= 5421) && (pixel_index <= 5465)) || ((pixel_index >= 5517) && (pixel_index <= 5561)) || ((pixel_index >= 5613) && (pixel_index <= 5657)) || ((pixel_index >= 5709) && (pixel_index <= 5753)) || ((pixel_index >= 5805) && (pixel_index <= 5849)) || ((pixel_index >= 5901) && (pixel_index <= 5945)) || ((pixel_index >= 5998) && (pixel_index <= 6041)) || (pixel_index >= 6094) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 25) begin
            if (((pixel_index >= 5) && (pixel_index <= 6)) || ((pixel_index >= 31) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 102)) || ((pixel_index >= 127) && (pixel_index <= 185)) || pixel_index == 197 || ((pixel_index >= 224) && (pixel_index <= 281)) || pixel_index == 293 || ((pixel_index >= 321) && (pixel_index <= 377)) || ((pixel_index >= 418) && (pixel_index <= 473)) || ((pixel_index >= 514) && (pixel_index <= 569)) || ((pixel_index >= 610) && (pixel_index <= 665)) || ((pixel_index >= 707) && (pixel_index <= 761)) || ((pixel_index >= 803) && (pixel_index <= 857)) || ((pixel_index >= 899) && (pixel_index <= 953)) || ((pixel_index >= 995) && (pixel_index <= 1049)) || ((pixel_index >= 1091) && (pixel_index <= 1145)) || ((pixel_index >= 1187) && (pixel_index <= 1241)) || ((pixel_index >= 1282) && (pixel_index <= 1337)) || ((pixel_index >= 1377) && (pixel_index <= 1433)) || ((pixel_index >= 1471) && (pixel_index <= 1529)) || ((pixel_index >= 1566) && (pixel_index <= 1625)) || ((pixel_index >= 1663) && (pixel_index <= 1721)) || ((pixel_index >= 1759) && (pixel_index <= 1817)) || ((pixel_index >= 1854) && (pixel_index <= 1913)) || ((pixel_index >= 1949) && (pixel_index <= 2009)) || ((pixel_index >= 2045) && (pixel_index <= 2105)) || ((pixel_index >= 2141) && (pixel_index <= 2201)) || ((pixel_index >= 2237) && (pixel_index <= 2297)) || ((pixel_index >= 2333) && (pixel_index <= 2393)) || ((pixel_index >= 2429) && (pixel_index <= 2489)) || pixel_index == 2502 || pixel_index == 2522 || ((pixel_index >= 2525) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2598)) || pixel_index == 2618 || ((pixel_index >= 2621) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2695)) || ((pixel_index >= 2717) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2792)) || ((pixel_index >= 2813) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2888)) || ((pixel_index >= 2909) && (pixel_index <= 2969)) || ((pixel_index >= 2981) && (pixel_index <= 2985)) || ((pixel_index >= 3005) && (pixel_index <= 3065)) || ((pixel_index >= 3077) && (pixel_index <= 3081)) || ((pixel_index >= 3101) && (pixel_index <= 3161)) || ((pixel_index >= 3173) && (pixel_index <= 3177)) || ((pixel_index >= 3199) && (pixel_index <= 3257)) || ((pixel_index >= 3269) && (pixel_index <= 3273)) || ((pixel_index >= 3295) && (pixel_index <= 3325)) || ((pixel_index >= 3327) && (pixel_index <= 3353)) || ((pixel_index >= 3365) && (pixel_index <= 3369)) || ((pixel_index >= 3391) && (pixel_index <= 3419)) || ((pixel_index >= 3426) && (pixel_index <= 3449)) || ((pixel_index >= 3461) && (pixel_index <= 3465)) || ((pixel_index >= 3488) && (pixel_index <= 3514)) || ((pixel_index >= 3523) && (pixel_index <= 3545)) || ((pixel_index >= 3557) && (pixel_index <= 3561)) || ((pixel_index >= 3585) && (pixel_index <= 3609)) || ((pixel_index >= 3620) && (pixel_index <= 3641)) || ((pixel_index >= 3653) && (pixel_index <= 3657)) || ((pixel_index >= 3682) && (pixel_index <= 3705)) || ((pixel_index >= 3716) && (pixel_index <= 3737)) || ((pixel_index >= 3749) && (pixel_index <= 3753)) || ((pixel_index >= 3780) && (pixel_index <= 3801)) || ((pixel_index >= 3812) && (pixel_index <= 3833)) || ((pixel_index >= 3845) && (pixel_index <= 3849)) || ((pixel_index >= 3877) && (pixel_index <= 3892)) || ((pixel_index >= 3895) && (pixel_index <= 3897)) || ((pixel_index >= 3908) && (pixel_index <= 3929)) || ((pixel_index >= 3941) && (pixel_index <= 3944)) || pixel_index == 3975 || pixel_index == 3992 || ((pixel_index >= 4004) && (pixel_index <= 4025)) || ((pixel_index >= 4037) && (pixel_index <= 4040)) || ((pixel_index >= 4100) && (pixel_index <= 4121)) || ((pixel_index >= 4133) && (pixel_index <= 4136)) || ((pixel_index >= 4195) && (pixel_index <= 4217)) || ((pixel_index >= 4229) && (pixel_index <= 4232)) || ((pixel_index >= 4291) && (pixel_index <= 4313)) || ((pixel_index >= 4325) && (pixel_index <= 4328)) || ((pixel_index >= 4386) && (pixel_index <= 4409)) || ((pixel_index >= 4421) && (pixel_index <= 4424)) || ((pixel_index >= 4480) && (pixel_index <= 4505)) || ((pixel_index >= 4517) && (pixel_index <= 4520)) || ((pixel_index >= 4570) && (pixel_index <= 4572)) || ((pixel_index >= 4575) && (pixel_index <= 4601)) || ((pixel_index >= 4613) && (pixel_index <= 4616)) || ((pixel_index >= 4666) && (pixel_index <= 4697)) || ((pixel_index >= 4709) && (pixel_index <= 4712)) || ((pixel_index >= 4762) && (pixel_index <= 4793)) || ((pixel_index >= 4805) && (pixel_index <= 4808)) || ((pixel_index >= 4858) && (pixel_index <= 4889)) || ((pixel_index >= 4901) && (pixel_index <= 4904)) || ((pixel_index >= 4954) && (pixel_index <= 4985)) || ((pixel_index >= 4997) && (pixel_index <= 5000)) || ((pixel_index >= 5050) && (pixel_index <= 5081)) || ((pixel_index >= 5093) && (pixel_index <= 5096)) || ((pixel_index >= 5146) && (pixel_index <= 5177)) || ((pixel_index >= 5189) && (pixel_index <= 5192)) || ((pixel_index >= 5242) && (pixel_index <= 5273)) || ((pixel_index >= 5285) && (pixel_index <= 5288)) || ((pixel_index >= 5338) && (pixel_index <= 5369)) || ((pixel_index >= 5381) && (pixel_index <= 5384)) || ((pixel_index >= 5434) && (pixel_index <= 5465)) || ((pixel_index >= 5477) && (pixel_index <= 5480)) || ((pixel_index >= 5530) && (pixel_index <= 5561)) || ((pixel_index >= 5573) && (pixel_index <= 5576)) || ((pixel_index >= 5626) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5671)) || ((pixel_index >= 5722) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5767)) || ((pixel_index >= 5817) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5863)) || ((pixel_index >= 5913) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 5959)) || ((pixel_index >= 6009) && (pixel_index <= 6041)) || ((pixel_index >= 6053) && (pixel_index <= 6055)) || (pixel_index >= 6105) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 26) begin
            if (((pixel_index >= 5) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 377)) || ((pixel_index >= 389) && (pixel_index <= 473)) || ((pixel_index >= 485) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 612)) || ((pixel_index >= 614) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 706)) || ((pixel_index >= 711) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 797)) || ((pixel_index >= 808) && (pixel_index <= 857)) || ((pixel_index >= 869) && (pixel_index <= 892)) || ((pixel_index >= 905) && (pixel_index <= 953)) || ((pixel_index >= 965) && (pixel_index <= 987)) || ((pixel_index >= 1002) && (pixel_index <= 1049)) || ((pixel_index >= 1061) && (pixel_index <= 1082)) || ((pixel_index >= 1098) && (pixel_index <= 1145)) || ((pixel_index >= 1157) && (pixel_index <= 1178)) || ((pixel_index >= 1195) && (pixel_index <= 1241)) || ((pixel_index >= 1253) && (pixel_index <= 1274)) || ((pixel_index >= 1292) && (pixel_index <= 1337)) || ((pixel_index >= 1349) && (pixel_index <= 1369)) || ((pixel_index >= 1389) && (pixel_index <= 1433)) || ((pixel_index >= 1445) && (pixel_index <= 1465)) || ((pixel_index >= 1486) && (pixel_index <= 1529)) || ((pixel_index >= 1541) && (pixel_index <= 1561)) || ((pixel_index >= 1582) && (pixel_index <= 1625)) || ((pixel_index >= 1637) && (pixel_index <= 1656)) || ((pixel_index >= 1678) && (pixel_index <= 1721)) || ((pixel_index >= 1733) && (pixel_index <= 1752)) || ((pixel_index >= 1774) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1848)) || ((pixel_index >= 1870) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 1944)) || ((pixel_index >= 1966) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2039)) || ((pixel_index >= 2062) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2135)) || ((pixel_index >= 2156) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2231)) || ((pixel_index >= 2251) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2327)) || ((pixel_index >= 2347) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2423)) || ((pixel_index >= 2443) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2519)) || ((pixel_index >= 2538) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2615)) || ((pixel_index >= 2633) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2711)) || ((pixel_index >= 2729) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2807)) || ((pixel_index >= 2825) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2903)) || ((pixel_index >= 2921) && (pixel_index <= 2969)) || ((pixel_index >= 2981) && (pixel_index <= 2999)) || ((pixel_index >= 3016) && (pixel_index <= 3065)) || ((pixel_index >= 3077) && (pixel_index <= 3095)) || ((pixel_index >= 3112) && (pixel_index <= 3161)) || ((pixel_index >= 3173) && (pixel_index <= 3194)) || ((pixel_index >= 3209) && (pixel_index <= 3230)) || ((pixel_index >= 3236) && (pixel_index <= 3257)) || ((pixel_index >= 3269) && (pixel_index <= 3291)) || ((pixel_index >= 3305) && (pixel_index <= 3326)) || ((pixel_index >= 3333) && (pixel_index <= 3353)) || ((pixel_index >= 3365) && (pixel_index <= 3388)) || ((pixel_index >= 3402) && (pixel_index <= 3421)) || ((pixel_index >= 3430) && (pixel_index <= 3449)) || ((pixel_index >= 3461) && (pixel_index <= 3484)) || ((pixel_index >= 3500) && (pixel_index <= 3517)) || ((pixel_index >= 3526) && (pixel_index <= 3545)) || ((pixel_index >= 3557) && (pixel_index <= 3581)) || ((pixel_index >= 3597) && (pixel_index <= 3613)) || ((pixel_index >= 3622) && (pixel_index <= 3641)) || ((pixel_index >= 3653) && (pixel_index <= 3677)) || ((pixel_index >= 3694) && (pixel_index <= 3710)) || ((pixel_index >= 3718) && (pixel_index <= 3737)) || ((pixel_index >= 3749) && (pixel_index <= 3773)) || ((pixel_index >= 3792) && (pixel_index <= 3801)) || ((pixel_index >= 3813) && (pixel_index <= 3833)) || ((pixel_index >= 3845) && (pixel_index <= 3868)) || ((pixel_index >= 3890) && (pixel_index <= 3891)) || ((pixel_index >= 3909) && (pixel_index <= 3929)) || ((pixel_index >= 3941) && (pixel_index <= 3965)) || ((pixel_index >= 4004) && (pixel_index <= 4025)) || ((pixel_index >= 4037) && (pixel_index <= 4061)) || ((pixel_index >= 4097) && (pixel_index <= 4121)) || ((pixel_index >= 4133) && (pixel_index <= 4157)) || ((pixel_index >= 4192) && (pixel_index <= 4217)) || ((pixel_index >= 4229) && (pixel_index <= 4253)) || ((pixel_index >= 4288) && (pixel_index <= 4313)) || ((pixel_index >= 4325) && (pixel_index <= 4349)) || ((pixel_index >= 4384) && (pixel_index <= 4409)) || ((pixel_index >= 4421) && (pixel_index <= 4445)) || ((pixel_index >= 4480) && (pixel_index <= 4505)) || ((pixel_index >= 4517) && (pixel_index <= 4541)) || ((pixel_index >= 4555) && (pixel_index <= 4556)) || ((pixel_index >= 4576) && (pixel_index <= 4601)) || ((pixel_index >= 4613) && (pixel_index <= 4637)) || ((pixel_index >= 4651) && (pixel_index <= 4652)) || ((pixel_index >= 4672) && (pixel_index <= 4697)) || ((pixel_index >= 4709) && (pixel_index <= 4733)) || ((pixel_index >= 4747) && (pixel_index <= 4748)) || ((pixel_index >= 4769) && (pixel_index <= 4793)) || ((pixel_index >= 4805) && (pixel_index <= 4829)) || ((pixel_index >= 4843) && (pixel_index <= 4844)) || ((pixel_index >= 4865) && (pixel_index <= 4889)) || ((pixel_index >= 4901) && (pixel_index <= 4925)) || pixel_index == 4940 || ((pixel_index >= 4960) && (pixel_index <= 4985)) || ((pixel_index >= 4997) && (pixel_index <= 5020)) || pixel_index == 5036 || ((pixel_index >= 5056) && (pixel_index <= 5081)) || ((pixel_index >= 5093) && (pixel_index <= 5116)) || pixel_index == 5132 || ((pixel_index >= 5152) && (pixel_index <= 5177)) || ((pixel_index >= 5189) && (pixel_index <= 5212)) || pixel_index == 5228 || ((pixel_index >= 5248) && (pixel_index <= 5273)) || ((pixel_index >= 5285) && (pixel_index <= 5308)) || ((pixel_index >= 5324) && (pixel_index <= 5325)) || ((pixel_index >= 5344) && (pixel_index <= 5369)) || ((pixel_index >= 5381) && (pixel_index <= 5404)) || ((pixel_index >= 5420) && (pixel_index <= 5421)) || ((pixel_index >= 5440) && (pixel_index <= 5465)) || ((pixel_index >= 5477) && (pixel_index <= 5500)) || ((pixel_index >= 5516) && (pixel_index <= 5517)) || ((pixel_index >= 5535) && (pixel_index <= 5561)) || ((pixel_index >= 5573) && (pixel_index <= 5595)) || ((pixel_index >= 5612) && (pixel_index <= 5613)) || ((pixel_index >= 5631) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5691)) || ((pixel_index >= 5707) && (pixel_index <= 5709)) || ((pixel_index >= 5727) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5787)) || ((pixel_index >= 5803) && (pixel_index <= 5805)) || ((pixel_index >= 5822) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5882)) || ((pixel_index >= 5898) && (pixel_index <= 5901)) || ((pixel_index >= 5917) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 5978)) || ((pixel_index >= 5994) && (pixel_index <= 5998)) || ((pixel_index >= 6012) && (pixel_index <= 6041)) || ((pixel_index >= 6053) && (pixel_index <= 6074)) || ((pixel_index >= 6090) && (pixel_index <= 6094)) || (pixel_index >= 6104) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 27) begin
            if (((pixel_index >= 5) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 377)) || ((pixel_index >= 389) && (pixel_index <= 473)) || ((pixel_index >= 485) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 857)) || ((pixel_index >= 869) && (pixel_index <= 902)) || ((pixel_index >= 906) && (pixel_index <= 953)) || ((pixel_index >= 965) && (pixel_index <= 992)) || ((pixel_index >= 1003) && (pixel_index <= 1049)) || ((pixel_index >= 1061) && (pixel_index <= 1087)) || ((pixel_index >= 1100) && (pixel_index <= 1145)) || ((pixel_index >= 1157) && (pixel_index <= 1182)) || ((pixel_index >= 1196) && (pixel_index <= 1241)) || ((pixel_index >= 1253) && (pixel_index <= 1278)) || ((pixel_index >= 1293) && (pixel_index <= 1337)) || ((pixel_index >= 1349) && (pixel_index <= 1373)) || ((pixel_index >= 1390) && (pixel_index <= 1433)) || ((pixel_index >= 1445) && (pixel_index <= 1469)) || ((pixel_index >= 1487) && (pixel_index <= 1529)) || ((pixel_index >= 1541) && (pixel_index <= 1565)) || ((pixel_index >= 1583) && (pixel_index <= 1625)) || ((pixel_index >= 1637) && (pixel_index <= 1660)) || ((pixel_index >= 1680) && (pixel_index <= 1721)) || ((pixel_index >= 1733) && (pixel_index <= 1756)) || ((pixel_index >= 1776) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1852)) || ((pixel_index >= 1872) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 1947)) || ((pixel_index >= 1968) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2043)) || ((pixel_index >= 2064) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2139)) || ((pixel_index >= 2160) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2235)) || ((pixel_index >= 2255) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2331)) || ((pixel_index >= 2349) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2427)) || ((pixel_index >= 2445) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2523)) || ((pixel_index >= 2541) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2619)) || ((pixel_index >= 2636) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2715)) || ((pixel_index >= 2731) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2810)) || ((pixel_index >= 2827) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2907)) || ((pixel_index >= 2923) && (pixel_index <= 2969)) || ((pixel_index >= 2981) && (pixel_index <= 3003)) || ((pixel_index >= 3019) && (pixel_index <= 3065)) || ((pixel_index >= 3077) && (pixel_index <= 3099)) || ((pixel_index >= 3114) && (pixel_index <= 3161)) || ((pixel_index >= 3173) && (pixel_index <= 3197)) || ((pixel_index >= 3210) && (pixel_index <= 3231)) || ((pixel_index >= 3234) && (pixel_index <= 3257)) || ((pixel_index >= 3269) && (pixel_index <= 3294)) || ((pixel_index >= 3307) && (pixel_index <= 3325)) || ((pixel_index >= 3332) && (pixel_index <= 3353)) || ((pixel_index >= 3365) && (pixel_index <= 3391)) || ((pixel_index >= 3403) && (pixel_index <= 3421)) || ((pixel_index >= 3429) && (pixel_index <= 3449)) || ((pixel_index >= 3461) && (pixel_index <= 3487)) || ((pixel_index >= 3500) && (pixel_index <= 3517)) || ((pixel_index >= 3525) && (pixel_index <= 3545)) || ((pixel_index >= 3557) && (pixel_index <= 3583)) || ((pixel_index >= 3598) && (pixel_index <= 3613)) || ((pixel_index >= 3621) && (pixel_index <= 3641)) || ((pixel_index >= 3653) && (pixel_index <= 3680)) || ((pixel_index >= 3695) && (pixel_index <= 3709)) || ((pixel_index >= 3717) && (pixel_index <= 3737)) || ((pixel_index >= 3749) && (pixel_index <= 3775)) || ((pixel_index >= 3792) && (pixel_index <= 3802)) || ((pixel_index >= 3813) && (pixel_index <= 3833)) || ((pixel_index >= 3845) && (pixel_index <= 3870)) || ((pixel_index >= 3889) && (pixel_index <= 3894)) || ((pixel_index >= 3908) && (pixel_index <= 3929)) || ((pixel_index >= 3941) && (pixel_index <= 3967)) || pixel_index == 3987 || ((pixel_index >= 4003) && (pixel_index <= 4025)) || ((pixel_index >= 4037) && (pixel_index <= 4064)) || ((pixel_index >= 4096) && (pixel_index <= 4121)) || ((pixel_index >= 4133) && (pixel_index <= 4160)) || ((pixel_index >= 4192) && (pixel_index <= 4217)) || ((pixel_index >= 4229) && (pixel_index <= 4255)) || ((pixel_index >= 4288) && (pixel_index <= 4313)) || ((pixel_index >= 4325) && (pixel_index <= 4351)) || ((pixel_index >= 4384) && (pixel_index <= 4409)) || ((pixel_index >= 4421) && (pixel_index <= 4447)) || pixel_index == 4461 || ((pixel_index >= 4481) && (pixel_index <= 4505)) || ((pixel_index >= 4517) && (pixel_index <= 4543)) || pixel_index == 4557 || ((pixel_index >= 4577) && (pixel_index <= 4601)) || ((pixel_index >= 4613) && (pixel_index <= 4639)) || ((pixel_index >= 4653) && (pixel_index <= 4654)) || ((pixel_index >= 4673) && (pixel_index <= 4697)) || ((pixel_index >= 4709) && (pixel_index <= 4735)) || ((pixel_index >= 4749) && (pixel_index <= 4750)) || ((pixel_index >= 4769) && (pixel_index <= 4793)) || ((pixel_index >= 4805) && (pixel_index <= 4831)) || ((pixel_index >= 4845) && (pixel_index <= 4846)) || ((pixel_index >= 4865) && (pixel_index <= 4889)) || ((pixel_index >= 4901) && (pixel_index <= 4926)) || ((pixel_index >= 4941) && (pixel_index <= 4943)) || ((pixel_index >= 4961) && (pixel_index <= 4985)) || ((pixel_index >= 4997) && (pixel_index <= 5022)) || ((pixel_index >= 5037) && (pixel_index <= 5039)) || ((pixel_index >= 5057) && (pixel_index <= 5081)) || ((pixel_index >= 5093) && (pixel_index <= 5118)) || ((pixel_index >= 5133) && (pixel_index <= 5135)) || ((pixel_index >= 5153) && (pixel_index <= 5177)) || ((pixel_index >= 5189) && (pixel_index <= 5214)) || ((pixel_index >= 5230) && (pixel_index <= 5231)) || ((pixel_index >= 5249) && (pixel_index <= 5273)) || ((pixel_index >= 5285) && (pixel_index <= 5310)) || ((pixel_index >= 5325) && (pixel_index <= 5327)) || ((pixel_index >= 5345) && (pixel_index <= 5369)) || ((pixel_index >= 5381) && (pixel_index <= 5406)) || ((pixel_index >= 5422) && (pixel_index <= 5423)) || ((pixel_index >= 5441) && (pixel_index <= 5465)) || ((pixel_index >= 5477) && (pixel_index <= 5502)) || ((pixel_index >= 5518) && (pixel_index <= 5520)) || ((pixel_index >= 5537) && (pixel_index <= 5561)) || ((pixel_index >= 5573) && (pixel_index <= 5598)) || ((pixel_index >= 5613) && (pixel_index <= 5616)) || ((pixel_index >= 5633) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5693)) || ((pixel_index >= 5709) && (pixel_index <= 5712)) || ((pixel_index >= 5729) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5789)) || ((pixel_index >= 5804) && (pixel_index <= 5808)) || ((pixel_index >= 5825) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5885)) || ((pixel_index >= 5900) && (pixel_index <= 5905)) || ((pixel_index >= 5920) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 5981)) || ((pixel_index >= 5996) && (pixel_index <= 6001)) || ((pixel_index >= 6015) && (pixel_index <= 6041)) || ((pixel_index >= 6053) && (pixel_index <= 6076)) || ((pixel_index >= 6092) && (pixel_index <= 6098)) || (pixel_index >= 6107) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 28) begin
            if (((pixel_index >= 5) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 377)) || ((pixel_index >= 389) && (pixel_index <= 473)) || ((pixel_index >= 485) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 857)) || ((pixel_index >= 869) && (pixel_index <= 953)) || ((pixel_index >= 965) && (pixel_index <= 1049)) || ((pixel_index >= 1061) && (pixel_index <= 1093)) || ((pixel_index >= 1095) && (pixel_index <= 1097)) || ((pixel_index >= 1100) && (pixel_index <= 1145)) || ((pixel_index >= 1157) && (pixel_index <= 1187)) || ((pixel_index >= 1198) && (pixel_index <= 1241)) || ((pixel_index >= 1253) && (pixel_index <= 1282)) || ((pixel_index >= 1295) && (pixel_index <= 1337)) || ((pixel_index >= 1349) && (pixel_index <= 1377)) || ((pixel_index >= 1392) && (pixel_index <= 1433)) || ((pixel_index >= 1445) && (pixel_index <= 1473)) || ((pixel_index >= 1488) && (pixel_index <= 1529)) || ((pixel_index >= 1541) && (pixel_index <= 1568)) || ((pixel_index >= 1584) && (pixel_index <= 1625)) || ((pixel_index >= 1637) && (pixel_index <= 1664)) || ((pixel_index >= 1681) && (pixel_index <= 1721)) || ((pixel_index >= 1733) && (pixel_index <= 1760)) || ((pixel_index >= 1778) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1855)) || ((pixel_index >= 1874) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 1951)) || ((pixel_index >= 1970) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2047)) || ((pixel_index >= 2066) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2142)) || ((pixel_index >= 2162) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2238)) || ((pixel_index >= 2258) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2334)) || ((pixel_index >= 2353) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2430)) || ((pixel_index >= 2448) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2526)) || ((pixel_index >= 2542) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2622)) || ((pixel_index >= 2639) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2718)) || ((pixel_index >= 2733) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2814)) || ((pixel_index >= 2829) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2910)) || pixel_index == 2921 || ((pixel_index >= 2925) && (pixel_index <= 2969)) || ((pixel_index >= 2981) && (pixel_index <= 3006)) || ((pixel_index >= 3021) && (pixel_index <= 3065)) || ((pixel_index >= 3077) && (pixel_index <= 3104)) || ((pixel_index >= 3117) && (pixel_index <= 3161)) || ((pixel_index >= 3173) && (pixel_index <= 3200)) || ((pixel_index >= 3213) && (pixel_index <= 3257)) || ((pixel_index >= 3269) && (pixel_index <= 3298)) || ((pixel_index >= 3309) && (pixel_index <= 3322)) || ((pixel_index >= 3327) && (pixel_index <= 3353)) || ((pixel_index >= 3365) && (pixel_index <= 3394)) || ((pixel_index >= 3405) && (pixel_index <= 3418)) || ((pixel_index >= 3424) && (pixel_index <= 3449)) || ((pixel_index >= 3461) && (pixel_index <= 3490)) || ((pixel_index >= 3502) && (pixel_index <= 3513)) || ((pixel_index >= 3521) && (pixel_index <= 3545)) || ((pixel_index >= 3557) && (pixel_index <= 3586)) || ((pixel_index >= 3598) && (pixel_index <= 3609)) || ((pixel_index >= 3617) && (pixel_index <= 3641)) || ((pixel_index >= 3653) && (pixel_index <= 3682)) || ((pixel_index >= 3695) && (pixel_index <= 3705)) || ((pixel_index >= 3713) && (pixel_index <= 3737)) || ((pixel_index >= 3749) && (pixel_index <= 3778)) || ((pixel_index >= 3791) && (pixel_index <= 3801)) || ((pixel_index >= 3809) && (pixel_index <= 3833)) || ((pixel_index >= 3845) && (pixel_index <= 3873)) || ((pixel_index >= 3888) && (pixel_index <= 3895)) || ((pixel_index >= 3904) && (pixel_index <= 3929)) || ((pixel_index >= 3941) && (pixel_index <= 3970)) || ((pixel_index >= 3984) && (pixel_index <= 3989)) || ((pixel_index >= 4000) && (pixel_index <= 4025)) || ((pixel_index >= 4037) && (pixel_index <= 4066)) || ((pixel_index >= 4081) && (pixel_index <= 4083)) || ((pixel_index >= 4093) && (pixel_index <= 4121)) || ((pixel_index >= 4133) && (pixel_index <= 4162)) || pixel_index == 4178 || ((pixel_index >= 4188) && (pixel_index <= 4217)) || ((pixel_index >= 4229) && (pixel_index <= 4258)) || ((pixel_index >= 4285) && (pixel_index <= 4313)) || ((pixel_index >= 4325) && (pixel_index <= 4354)) || ((pixel_index >= 4381) && (pixel_index <= 4409)) || ((pixel_index >= 4421) && (pixel_index <= 4450)) || ((pixel_index >= 4478) && (pixel_index <= 4505)) || ((pixel_index >= 4517) && (pixel_index <= 4546)) || ((pixel_index >= 4574) && (pixel_index <= 4601)) || ((pixel_index >= 4613) && (pixel_index <= 4642)) || ((pixel_index >= 4671) && (pixel_index <= 4697)) || ((pixel_index >= 4709) && (pixel_index <= 4738)) || ((pixel_index >= 4767) && (pixel_index <= 4793)) || ((pixel_index >= 4805) && (pixel_index <= 4833)) || ((pixel_index >= 4863) && (pixel_index <= 4889)) || ((pixel_index >= 4901) && (pixel_index <= 4929)) || ((pixel_index >= 4960) && (pixel_index <= 4985)) || ((pixel_index >= 4997) && (pixel_index <= 5025)) || ((pixel_index >= 5056) && (pixel_index <= 5081)) || ((pixel_index >= 5093) && (pixel_index <= 5121)) || ((pixel_index >= 5152) && (pixel_index <= 5177)) || ((pixel_index >= 5189) && (pixel_index <= 5217)) || ((pixel_index >= 5249) && (pixel_index <= 5273)) || ((pixel_index >= 5285) && (pixel_index <= 5313)) || ((pixel_index >= 5345) && (pixel_index <= 5369)) || ((pixel_index >= 5381) && (pixel_index <= 5409)) || pixel_index == 5423 || ((pixel_index >= 5441) && (pixel_index <= 5465)) || ((pixel_index >= 5477) && (pixel_index <= 5505)) || pixel_index == 5519 || ((pixel_index >= 5537) && (pixel_index <= 5561)) || ((pixel_index >= 5573) && (pixel_index <= 5600)) || ((pixel_index >= 5614) && (pixel_index <= 5616)) || ((pixel_index >= 5633) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5696)) || ((pixel_index >= 5710) && (pixel_index <= 5712)) || ((pixel_index >= 5729) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5792)) || ((pixel_index >= 5806) && (pixel_index <= 5808)) || ((pixel_index >= 5825) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5887)) || ((pixel_index >= 5902) && (pixel_index <= 5905)) || ((pixel_index >= 5920) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 5983)) || ((pixel_index >= 5999) && (pixel_index <= 6001)) || ((pixel_index >= 6013) && (pixel_index <= 6041)) || ((pixel_index >= 6053) && (pixel_index <= 6079)) || ((pixel_index >= 6095) && (pixel_index <= 6098)) || (pixel_index >= 6108) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 29) begin
            if (((pixel_index >= 5) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 377)) || ((pixel_index >= 389) && (pixel_index <= 473)) || ((pixel_index >= 485) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 857)) || ((pixel_index >= 869) && (pixel_index <= 953)) || ((pixel_index >= 965) && (pixel_index <= 1049)) || ((pixel_index >= 1061) && (pixel_index <= 1093)) || ((pixel_index >= 1098) && (pixel_index <= 1145)) || ((pixel_index >= 1157) && (pixel_index <= 1188)) || pixel_index == 1198 || ((pixel_index >= 1206) && (pixel_index <= 1241)) || ((pixel_index >= 1253) && (pixel_index <= 1283)) || ((pixel_index >= 1303) && (pixel_index <= 1337)) || ((pixel_index >= 1349) && (pixel_index <= 1379)) || ((pixel_index >= 1399) && (pixel_index <= 1433)) || ((pixel_index >= 1445) && (pixel_index <= 1474)) || ((pixel_index >= 1494) && (pixel_index <= 1529)) || ((pixel_index >= 1541) && (pixel_index <= 1569)) || ((pixel_index >= 1590) && (pixel_index <= 1625)) || ((pixel_index >= 1637) && (pixel_index <= 1665)) || ((pixel_index >= 1685) && (pixel_index <= 1721)) || ((pixel_index >= 1733) && (pixel_index <= 1761)) || ((pixel_index >= 1780) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1857)) || ((pixel_index >= 1876) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 1951)) || ((pixel_index >= 1973) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2047)) || ((pixel_index >= 2069) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2144)) || ((pixel_index >= 2165) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2240)) || ((pixel_index >= 2260) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2336)) || ((pixel_index >= 2356) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2432)) || ((pixel_index >= 2451) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2528)) || ((pixel_index >= 2546) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2624)) || ((pixel_index >= 2642) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2719)) || ((pixel_index >= 2738) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2815)) || ((pixel_index >= 2834) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2912)) || ((pixel_index >= 2926) && (pixel_index <= 2927)) || ((pixel_index >= 2930) && (pixel_index <= 2969)) || ((pixel_index >= 2981) && (pixel_index <= 3008)) || ((pixel_index >= 3022) && (pixel_index <= 3023)) || ((pixel_index >= 3026) && (pixel_index <= 3065)) || ((pixel_index >= 3077) && (pixel_index <= 3108)) || pixel_index == 3119 || ((pixel_index >= 3121) && (pixel_index <= 3161)) || ((pixel_index >= 3173) && (pixel_index <= 3204)) || ((pixel_index >= 3217) && (pixel_index <= 3257)) || ((pixel_index >= 3269) && (pixel_index <= 3300)) || ((pixel_index >= 3313) && (pixel_index <= 3320)) || ((pixel_index >= 3324) && (pixel_index <= 3353)) || ((pixel_index >= 3365) && (pixel_index <= 3397)) || ((pixel_index >= 3409) && (pixel_index <= 3415)) || ((pixel_index >= 3421) && (pixel_index <= 3449)) || ((pixel_index >= 3461) && (pixel_index <= 3493)) || ((pixel_index >= 3506) && (pixel_index <= 3510)) || ((pixel_index >= 3517) && (pixel_index <= 3545)) || ((pixel_index >= 3557) && (pixel_index <= 3589)) || ((pixel_index >= 3602) && (pixel_index <= 3606)) || ((pixel_index >= 3614) && (pixel_index <= 3641)) || ((pixel_index >= 3653) && (pixel_index <= 3685)) || ((pixel_index >= 3699) && (pixel_index <= 3702)) || ((pixel_index >= 3710) && (pixel_index <= 3737)) || ((pixel_index >= 3749) && (pixel_index <= 3781)) || ((pixel_index >= 3795) && (pixel_index <= 3798)) || ((pixel_index >= 3805) && (pixel_index <= 3833)) || ((pixel_index >= 3845) && (pixel_index <= 3876)) || ((pixel_index >= 3891) && (pixel_index <= 3893)) || ((pixel_index >= 3901) && (pixel_index <= 3929)) || ((pixel_index >= 3941) && (pixel_index <= 3973)) || pixel_index == 3988 || ((pixel_index >= 3996) && (pixel_index <= 4025)) || ((pixel_index >= 4037) && (pixel_index <= 4069)) || ((pixel_index >= 4090) && (pixel_index <= 4121)) || ((pixel_index >= 4133) && (pixel_index <= 4165)) || ((pixel_index >= 4186) && (pixel_index <= 4217)) || ((pixel_index >= 4229) && (pixel_index <= 4261)) || ((pixel_index >= 4282) && (pixel_index <= 4313)) || ((pixel_index >= 4325) && (pixel_index <= 4357)) || ((pixel_index >= 4379) && (pixel_index <= 4409)) || ((pixel_index >= 4421) && (pixel_index <= 4452)) || ((pixel_index >= 4475) && (pixel_index <= 4505)) || ((pixel_index >= 4517) && (pixel_index <= 4548)) || ((pixel_index >= 4572) && (pixel_index <= 4601)) || ((pixel_index >= 4613) && (pixel_index <= 4644)) || ((pixel_index >= 4668) && (pixel_index <= 4697)) || ((pixel_index >= 4709) && (pixel_index <= 4740)) || ((pixel_index >= 4765) && (pixel_index <= 4793)) || ((pixel_index >= 4805) && (pixel_index <= 4836)) || ((pixel_index >= 4861) && (pixel_index <= 4889)) || ((pixel_index >= 4901) && (pixel_index <= 4932)) || ((pixel_index >= 4957) && (pixel_index <= 4985)) || ((pixel_index >= 4997) && (pixel_index <= 5028)) || ((pixel_index >= 5054) && (pixel_index <= 5081)) || ((pixel_index >= 5093) && (pixel_index <= 5124)) || ((pixel_index >= 5150) && (pixel_index <= 5177)) || ((pixel_index >= 5189) && (pixel_index <= 5219)) || ((pixel_index >= 5246) && (pixel_index <= 5273)) || ((pixel_index >= 5285) && (pixel_index <= 5315)) || ((pixel_index >= 5342) && (pixel_index <= 5369)) || ((pixel_index >= 5381) && (pixel_index <= 5411)) || ((pixel_index >= 5439) && (pixel_index <= 5465)) || ((pixel_index >= 5477) && (pixel_index <= 5508)) || ((pixel_index >= 5535) && (pixel_index <= 5561)) || ((pixel_index >= 5573) && (pixel_index <= 5604)) || ((pixel_index >= 5631) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5699)) || ((pixel_index >= 5727) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5795)) || ((pixel_index >= 5823) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5891)) || ((pixel_index >= 5918) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 5987)) || ((pixel_index >= 6013) && (pixel_index <= 6041)) || ((pixel_index >= 6053) && (pixel_index <= 6082)) || (pixel_index >= 6108) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 30) begin
            if (((pixel_index >= 5) && (pixel_index <= 34)) || ((pixel_index >= 41) && (pixel_index <= 89)) || ((pixel_index >= 101) && (pixel_index <= 129)) || ((pixel_index >= 138) && (pixel_index <= 185)) || ((pixel_index >= 197) && (pixel_index <= 225)) || ((pixel_index >= 235) && (pixel_index <= 281)) || ((pixel_index >= 293) && (pixel_index <= 320)) || ((pixel_index >= 336) && (pixel_index <= 337)) || ((pixel_index >= 349) && (pixel_index <= 377)) || ((pixel_index >= 389) && (pixel_index <= 416)) || ((pixel_index >= 445) && (pixel_index <= 473)) || ((pixel_index >= 485) && (pixel_index <= 511)) || ((pixel_index >= 541) && (pixel_index <= 569)) || ((pixel_index >= 581) && (pixel_index <= 607)) || ((pixel_index >= 637) && (pixel_index <= 665)) || ((pixel_index >= 677) && (pixel_index <= 702)) || ((pixel_index >= 733) && (pixel_index <= 761)) || ((pixel_index >= 773) && (pixel_index <= 798)) || ((pixel_index >= 829) && (pixel_index <= 857)) || ((pixel_index >= 869) && (pixel_index <= 894)) || ((pixel_index >= 924) && (pixel_index <= 953)) || ((pixel_index >= 965) && (pixel_index <= 989)) || ((pixel_index >= 1020) && (pixel_index <= 1049)) || ((pixel_index >= 1061) && (pixel_index <= 1085)) || ((pixel_index >= 1115) && (pixel_index <= 1145)) || ((pixel_index >= 1157) && (pixel_index <= 1182)) || ((pixel_index >= 1210) && (pixel_index <= 1241)) || ((pixel_index >= 1253) && (pixel_index <= 1279)) || ((pixel_index >= 1306) && (pixel_index <= 1337)) || ((pixel_index >= 1349) && (pixel_index <= 1374)) || ((pixel_index >= 1401) && (pixel_index <= 1433)) || ((pixel_index >= 1445) && (pixel_index <= 1469)) || ((pixel_index >= 1498) && (pixel_index <= 1529)) || ((pixel_index >= 1541) && (pixel_index <= 1564)) || ((pixel_index >= 1594) && (pixel_index <= 1625)) || ((pixel_index >= 1637) && (pixel_index <= 1660)) || ((pixel_index >= 1690) && (pixel_index <= 1721)) || ((pixel_index >= 1733) && (pixel_index <= 1758)) || ((pixel_index >= 1786) && (pixel_index <= 1817)) || ((pixel_index >= 1829) && (pixel_index <= 1855)) || ((pixel_index >= 1881) && (pixel_index <= 1913)) || ((pixel_index >= 1925) && (pixel_index <= 1951)) || ((pixel_index >= 1977) && (pixel_index <= 2009)) || ((pixel_index >= 2021) && (pixel_index <= 2047)) || ((pixel_index >= 2072) && (pixel_index <= 2105)) || ((pixel_index >= 2117) && (pixel_index <= 2143)) || ((pixel_index >= 2167) && (pixel_index <= 2201)) || ((pixel_index >= 2213) && (pixel_index <= 2239)) || ((pixel_index >= 2262) && (pixel_index <= 2297)) || ((pixel_index >= 2309) && (pixel_index <= 2334)) || ((pixel_index >= 2358) && (pixel_index <= 2393)) || ((pixel_index >= 2405) && (pixel_index <= 2430)) || ((pixel_index >= 2455) && (pixel_index <= 2489)) || ((pixel_index >= 2501) && (pixel_index <= 2527)) || ((pixel_index >= 2551) && (pixel_index <= 2585)) || ((pixel_index >= 2597) && (pixel_index <= 2623)) || pixel_index == 2643 || ((pixel_index >= 2647) && (pixel_index <= 2681)) || ((pixel_index >= 2693) && (pixel_index <= 2719)) || pixel_index == 2739 || ((pixel_index >= 2743) && (pixel_index <= 2777)) || ((pixel_index >= 2789) && (pixel_index <= 2815)) || ((pixel_index >= 2834) && (pixel_index <= 2835)) || ((pixel_index >= 2839) && (pixel_index <= 2873)) || ((pixel_index >= 2885) && (pixel_index <= 2911)) || pixel_index == 2915 || ((pixel_index >= 2930) && (pixel_index <= 2931)) || ((pixel_index >= 2935) && (pixel_index <= 2969)) || ((pixel_index >= 2981) && (pixel_index <= 3011)) || pixel_index == 3027 || ((pixel_index >= 3031) && (pixel_index <= 3065)) || ((pixel_index >= 3077) && (pixel_index <= 3107)) || ((pixel_index >= 3123) && (pixel_index <= 3124)) || ((pixel_index >= 3127) && (pixel_index <= 3161)) || ((pixel_index >= 3173) && (pixel_index <= 3203)) || pixel_index == 3220 || ((pixel_index >= 3223) && (pixel_index <= 3257)) || ((pixel_index >= 3269) && (pixel_index <= 3299)) || ((pixel_index >= 3319) && (pixel_index <= 3353)) || ((pixel_index >= 3365) && (pixel_index <= 3394)) || ((pixel_index >= 3415) && (pixel_index <= 3417)) || ((pixel_index >= 3424) && (pixel_index <= 3449)) || ((pixel_index >= 3461) && (pixel_index <= 3490)) || ((pixel_index >= 3511) && (pixel_index <= 3512)) || ((pixel_index >= 3522) && (pixel_index <= 3545)) || ((pixel_index >= 3557) && (pixel_index <= 3587)) || ((pixel_index >= 3607) && (pixel_index <= 3608)) || ((pixel_index >= 3618) && (pixel_index <= 3641)) || ((pixel_index >= 3653) && (pixel_index <= 3683)) || ((pixel_index >= 3703) && (pixel_index <= 3704)) || ((pixel_index >= 3714) && (pixel_index <= 3737)) || ((pixel_index >= 3749) && (pixel_index <= 3779)) || ((pixel_index >= 3799) && (pixel_index <= 3800)) || ((pixel_index >= 3811) && (pixel_index <= 3833)) || ((pixel_index >= 3845) && (pixel_index <= 3875)) || pixel_index == 3896 || ((pixel_index >= 3906) && (pixel_index <= 3929)) || ((pixel_index >= 3941) && (pixel_index <= 3971)) || ((pixel_index >= 4002) && (pixel_index <= 4025)) || ((pixel_index >= 4037) && (pixel_index <= 4067)) || ((pixel_index >= 4098) && (pixel_index <= 4121)) || ((pixel_index >= 4133) && (pixel_index <= 4163)) || ((pixel_index >= 4193) && (pixel_index <= 4217)) || ((pixel_index >= 4229) && (pixel_index <= 4259)) || ((pixel_index >= 4289) && (pixel_index <= 4313)) || ((pixel_index >= 4325) && (pixel_index <= 4355)) || ((pixel_index >= 4384) && (pixel_index <= 4409)) || ((pixel_index >= 4421) && (pixel_index <= 4451)) || ((pixel_index >= 4476) && (pixel_index <= 4505)) || ((pixel_index >= 4517) && (pixel_index <= 4547)) || pixel_index == 4549 || ((pixel_index >= 4571) && (pixel_index <= 4601)) || ((pixel_index >= 4613) && (pixel_index <= 4643)) || ((pixel_index >= 4645) && (pixel_index <= 4646)) || ((pixel_index >= 4668) && (pixel_index <= 4697)) || ((pixel_index >= 4709) && (pixel_index <= 4739)) || ((pixel_index >= 4741) && (pixel_index <= 4742)) || ((pixel_index >= 4764) && (pixel_index <= 4793)) || ((pixel_index >= 4805) && (pixel_index <= 4835)) || ((pixel_index >= 4861) && (pixel_index <= 4889)) || ((pixel_index >= 4901) && (pixel_index <= 4930)) || ((pixel_index >= 4957) && (pixel_index <= 4985)) || ((pixel_index >= 4997) && (pixel_index <= 5027)) || pixel_index == 5029 || ((pixel_index >= 5053) && (pixel_index <= 5081)) || ((pixel_index >= 5093) && (pixel_index <= 5123)) || pixel_index == 5125 || ((pixel_index >= 5150) && (pixel_index <= 5177)) || ((pixel_index >= 5189) && (pixel_index <= 5219)) || ((pixel_index >= 5246) && (pixel_index <= 5273)) || ((pixel_index >= 5285) && (pixel_index <= 5315)) || ((pixel_index >= 5342) && (pixel_index <= 5369)) || ((pixel_index >= 5381) && (pixel_index <= 5411)) || ((pixel_index >= 5438) && (pixel_index <= 5465)) || ((pixel_index >= 5477) && (pixel_index <= 5507)) || ((pixel_index >= 5534) && (pixel_index <= 5561)) || ((pixel_index >= 5573) && (pixel_index <= 5603)) || ((pixel_index >= 5630) && (pixel_index <= 5657)) || ((pixel_index >= 5669) && (pixel_index <= 5699)) || ((pixel_index >= 5727) && (pixel_index <= 5753)) || ((pixel_index >= 5765) && (pixel_index <= 5795)) || ((pixel_index >= 5823) && (pixel_index <= 5849)) || ((pixel_index >= 5861) && (pixel_index <= 5891)) || ((pixel_index >= 5919) && (pixel_index <= 5945)) || ((pixel_index >= 5957) && (pixel_index <= 5987)) || ((pixel_index >= 6015) && (pixel_index <= 6041)) || ((pixel_index >= 6053) && (pixel_index <= 6083)) || (pixel_index >= 6111) && (pixel_index <= 6137)) oled_data = 16'b1111111111111111;
            else oled_data = 0;
        end
        else if (frame_count == 31) begin
            oled_data = 0;
            done = 1;
        end
    end
    
endmodule