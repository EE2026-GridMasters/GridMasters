`timescale 1ns / 1ps

module display_start(
    input [12:0] pixel_index,
    output reg [15:0] oled_data
    );
    
    parameter PINK_HEX = 16'hF899;
    parameter BG_BLUE_HEX = 16'b0000000001000100;
    
    always @(*) begin
        if ((pixel_index >= 208 && pixel_index <= 214) || (pixel_index >= 223 && pixel_index <= 225) || (pixel_index >= 240 && pixel_index <= 242) || (pixel_index >= 250 && pixel_index <= 256) || (pixel_index >= 264 && pixel_index <= 266) || (pixel_index >= 274 && pixel_index <= 276) || (pixel_index >= 304 && pixel_index <= 310) || (pixel_index >= 319 && pixel_index <= 321) || (pixel_index >= 336 && pixel_index <= 338) || (pixel_index >= 346 && pixel_index <= 352) || (pixel_index >= 360 && pixel_index <= 362) || (pixel_index >= 370 && pixel_index <= 372) || (pixel_index >= 400 && pixel_index <= 406) || (pixel_index >= 415 && pixel_index <= 417) || (pixel_index >= 432 && pixel_index <= 434) || (pixel_index >= 442 && pixel_index <= 448) || (pixel_index >= 456 && pixel_index <= 458) || (pixel_index >= 466 && pixel_index <= 468) || (pixel_index >= 493 && pixel_index <= 495) || (pixel_index >= 503 && pixel_index <= 505) || (pixel_index >= 511 && pixel_index <= 513) || (pixel_index >= 528 && pixel_index <= 530) || (pixel_index >= 535 && pixel_index <= 537) || (pixel_index >= 545 && pixel_index <= 547) || (pixel_index >= 552 && pixel_index <= 554) || (pixel_index >= 562 && pixel_index <= 564) || (pixel_index >= 589 && pixel_index <= 591) || (pixel_index >= 599 && pixel_index <= 601) || (pixel_index >= 607 && pixel_index <= 609) || (pixel_index >= 624 && pixel_index <= 626) || (pixel_index >= 631 && pixel_index <= 633) || (pixel_index >= 641 && pixel_index <= 643) || (pixel_index >= 648 && pixel_index <= 650) || (pixel_index >= 655 && pixel_index <= 657) || (pixel_index >= 685 && pixel_index <= 687) || (pixel_index >= 695 && pixel_index <= 697) || (pixel_index >= 703 && pixel_index <= 705) || (pixel_index >= 720 && pixel_index <= 722) || (pixel_index >= 727 && pixel_index <= 729) || (pixel_index >= 737 && pixel_index <= 739) || (pixel_index >= 744 && pixel_index <= 746) || (pixel_index >= 751 && pixel_index <= 753) || (pixel_index >= 781 && pixel_index <= 783) || (pixel_index >= 799 && pixel_index <= 801) || (pixel_index >= 816 && pixel_index <= 818) || (pixel_index >= 823 && pixel_index <= 825) || (pixel_index >= 840 && pixel_index <= 842) || (pixel_index >= 847 && pixel_index <= 849) || (pixel_index >= 877 && pixel_index <= 879) || (pixel_index >= 895 && pixel_index <= 897) || (pixel_index >= 912 && pixel_index <= 914) || (pixel_index >= 919 && pixel_index <= 921) || (pixel_index >= 936 && pixel_index <= 938) || (pixel_index >= 943 && pixel_index <= 945) || (pixel_index >= 973 && pixel_index <= 975) || (pixel_index >= 991 && pixel_index <= 993) || (pixel_index >= 1008 && pixel_index <= 1010) || (pixel_index >= 1015 && pixel_index <= 1017) || (pixel_index >= 1032 && pixel_index <= 1038) || (pixel_index >= 1069 && pixel_index <= 1071) || (pixel_index >= 1087 && pixel_index <= 1089) || (pixel_index >= 1104 && pixel_index <= 1106) || (pixel_index >= 1111 && pixel_index <= 1113) || (pixel_index >= 1128 && pixel_index <= 1134) || (pixel_index >= 1165 && pixel_index <= 1167) || (pixel_index >= 1183 && pixel_index <= 1185) || (pixel_index >= 1200 && pixel_index <= 1202) || (pixel_index >= 1207 && pixel_index <= 1209) || (pixel_index >= 1224 && pixel_index <= 1230) || (pixel_index >= 1261 && pixel_index <= 1263) || (pixel_index >= 1279 && pixel_index <= 1281) || (pixel_index >= 1296 && pixel_index <= 1298) || (pixel_index >= 1303 && pixel_index <= 1305) || (pixel_index >= 1320 && pixel_index <= 1322) || (pixel_index >= 1327 && pixel_index <= 1329) || (pixel_index >= 1357 && pixel_index <= 1359) || (pixel_index >= 1367 && pixel_index <= 1369) || (pixel_index >= 1375 && pixel_index <= 1377) || (pixel_index >= 1392 && pixel_index <= 1394) || (pixel_index >= 1399 && pixel_index <= 1401) || (pixel_index >= 1409 && pixel_index <= 1411) || (pixel_index >= 1416 && pixel_index <= 1418) || (pixel_index >= 1423 && pixel_index <= 1425) || (pixel_index >= 1453 && pixel_index <= 1455) || (pixel_index >= 1463 && pixel_index <= 1465) || (pixel_index >= 1471 && pixel_index <= 1473) || (pixel_index >= 1488 && pixel_index <= 1490) || (pixel_index >= 1495 && pixel_index <= 1497) || (pixel_index >= 1505 && pixel_index <= 1507) || (pixel_index >= 1512 && pixel_index <= 1514) || (pixel_index >= 1519 && pixel_index <= 1521) || (pixel_index >= 1549 && pixel_index <= 1551) || (pixel_index >= 1559 && pixel_index <= 1561) || (pixel_index >= 1567 && pixel_index <= 1569) || (pixel_index >= 1584 && pixel_index <= 1586) || (pixel_index >= 1591 && pixel_index <= 1593) || (pixel_index >= 1601 && pixel_index <= 1603) || (pixel_index >= 1608 && pixel_index <= 1610) || (pixel_index >= 1618 && pixel_index <= 1620) || (pixel_index >= 1648 && pixel_index <= 1654) || (pixel_index >= 1663 && pixel_index <= 1674) || (pixel_index >= 1680 && pixel_index <= 1682) || (pixel_index >= 1690 && pixel_index <= 1696) || (pixel_index >= 1704 && pixel_index <= 1706) || (pixel_index >= 1714 && pixel_index <= 1716) || (pixel_index >= 1744 && pixel_index <= 1750) || (pixel_index >= 1759 && pixel_index <= 1770) || (pixel_index >= 1776 && pixel_index <= 1778) || (pixel_index >= 1786 && pixel_index <= 1792) || (pixel_index >= 1800 && pixel_index <= 1802) || (pixel_index >= 1810 && pixel_index <= 1812) || (pixel_index >= 1840 && pixel_index <= 1846) || (pixel_index >= 1855 && pixel_index <= 1866) || (pixel_index >= 1872 && pixel_index <= 1874) || (pixel_index >= 1882 && pixel_index <= 1888) || (pixel_index >= 1896 && pixel_index <= 1898) || (pixel_index >= 1906 && pixel_index <= 1908) || (pixel_index >= 2242 && pixel_index <= 2254) || (pixel_index >= 2262 && pixel_index <= 2268) || (pixel_index >= 2338 && pixel_index <= 2350) || (pixel_index >= 2358 && pixel_index <= 2364) || (pixel_index >= 2434 && pixel_index <= 2446) || (pixel_index >= 2454 && pixel_index <= 2460) || (pixel_index >= 2535 && pixel_index <= 2537) || (pixel_index >= 2547 && pixel_index <= 2549) || (pixel_index >= 2557 && pixel_index <= 2559) || (pixel_index >= 2631 && pixel_index <= 2633) || (pixel_index >= 2643 && pixel_index <= 2645) || (pixel_index >= 2653 && pixel_index <= 2655) || (pixel_index >= 2727 && pixel_index <= 2729) || (pixel_index >= 2739 && pixel_index <= 2741) || (pixel_index >= 2749 && pixel_index <= 2751) || (pixel_index >= 2823 && pixel_index <= 2825) || (pixel_index >= 2835 && pixel_index <= 2837) || (pixel_index >= 2845 && pixel_index <= 2847) || (pixel_index >= 2919 && pixel_index <= 2921) || (pixel_index >= 2931 && pixel_index <= 2933) || (pixel_index >= 2941 && pixel_index <= 2943) || (pixel_index >= 3015 && pixel_index <= 3017) || (pixel_index >= 3027 && pixel_index <= 3029) || (pixel_index >= 3037 && pixel_index <= 3039) || (pixel_index >= 3111 && pixel_index <= 3113) || (pixel_index >= 3123 && pixel_index <= 3125) || (pixel_index >= 3133 && pixel_index <= 3135) || (pixel_index >= 3207 && pixel_index <= 3209) || (pixel_index >= 3219 && pixel_index <= 3221) || (pixel_index >= 3229 && pixel_index <= 3231) || (pixel_index >= 3303 && pixel_index <= 3305) || (pixel_index >= 3315 && pixel_index <= 3317) || (pixel_index >= 3325 && pixel_index <= 3327) || (pixel_index >= 3399 && pixel_index <= 3401) || (pixel_index >= 3411 && pixel_index <= 3413) || (pixel_index >= 3421 && pixel_index <= 3423) || (pixel_index >= 3495 && pixel_index <= 3497) || (pixel_index >= 3507 && pixel_index <= 3509) || (pixel_index >= 3517 && pixel_index <= 3519) || (pixel_index >= 3591 && pixel_index <= 3593) || (pixel_index >= 3603 && pixel_index <= 3605) || (pixel_index >= 3613 && pixel_index <= 3615) || (pixel_index >= 3687 && pixel_index <= 3689) || (pixel_index >= 3702 && pixel_index <= 3708) || (pixel_index >= 3783 && pixel_index <= 3785) || (pixel_index >= 3798 && pixel_index <= 3804) || (pixel_index >= 3879 && pixel_index <= 3881) || (pixel_index >= 3894 && pixel_index <= 3900) || (pixel_index >= 4232 && pixel_index <= 4238) || (pixel_index >= 4246 && pixel_index <= 4258) || (pixel_index >= 4266 && pixel_index <= 4272) || (pixel_index >= 4280 && pixel_index <= 4289) || (pixel_index >= 4297 && pixel_index <= 4309) || (pixel_index >= 4314 && pixel_index <= 4316) || (pixel_index >= 4328 && pixel_index <= 4334) || (pixel_index >= 4342 && pixel_index <= 4354) || (pixel_index >= 4362 && pixel_index <= 4368) || (pixel_index >= 4376 && pixel_index <= 4385) || (pixel_index >= 4393 && pixel_index <= 4405) || (pixel_index >= 4410 && pixel_index <= 4412) || (pixel_index >= 4424 && pixel_index <= 4430) || (pixel_index >= 4438 && pixel_index <= 4450) || (pixel_index >= 4458 && pixel_index <= 4464) || (pixel_index >= 4472 && pixel_index <= 4481) || (pixel_index >= 4489 && pixel_index <= 4501) || (pixel_index >= 4506 && pixel_index <= 4508) || (pixel_index >= 4517 && pixel_index <= 4519) || (pixel_index >= 4527 && pixel_index <= 4529) || (pixel_index >= 4539 && pixel_index <= 4541) || (pixel_index >= 4551 && pixel_index <= 4553) || (pixel_index >= 4561 && pixel_index <= 4563) || (pixel_index >= 4568 && pixel_index <= 4570) || (pixel_index >= 4578 && pixel_index <= 4580) || (pixel_index >= 4590 && pixel_index <= 4592) || (pixel_index >= 4602 && pixel_index <= 4604) || (pixel_index >= 4613 && pixel_index <= 4615) || (pixel_index >= 4623 && pixel_index <= 4625) || (pixel_index >= 4635 && pixel_index <= 4637) || (pixel_index >= 4647 && pixel_index <= 4649) || (pixel_index >= 4657 && pixel_index <= 4659) || (pixel_index >= 4664 && pixel_index <= 4666) || (pixel_index >= 4674 && pixel_index <= 4676) || (pixel_index >= 4686 && pixel_index <= 4688) || (pixel_index >= 4698 && pixel_index <= 4700) || (pixel_index >= 4709 && pixel_index <= 4711) || (pixel_index >= 4719 && pixel_index <= 4721) || (pixel_index >= 4731 && pixel_index <= 4733) || (pixel_index >= 4743 && pixel_index <= 4745) || (pixel_index >= 4753 && pixel_index <= 4755) || (pixel_index >= 4760 && pixel_index <= 4762) || (pixel_index >= 4770 && pixel_index <= 4772) || (pixel_index >= 4782 && pixel_index <= 4784) || (pixel_index >= 4794 && pixel_index <= 4796) || (pixel_index >= 4805 && pixel_index <= 4807) || (pixel_index >= 4815 && pixel_index <= 4817) || (pixel_index >= 4827 && pixel_index <= 4829) || (pixel_index >= 4839 && pixel_index <= 4841) || (pixel_index >= 4849 && pixel_index <= 4851) || (pixel_index >= 4856 && pixel_index <= 4858) || (pixel_index >= 4866 && pixel_index <= 4868) || (pixel_index >= 4878 && pixel_index <= 4880) || (pixel_index >= 4890 && pixel_index <= 4892) || (pixel_index >= 4901 && pixel_index <= 4903) || (pixel_index >= 4923 && pixel_index <= 4925) || (pixel_index >= 4935 && pixel_index <= 4937) || (pixel_index >= 4945 && pixel_index <= 4947) || (pixel_index >= 4952 && pixel_index <= 4954) || (pixel_index >= 4962 && pixel_index <= 4964) || (pixel_index >= 4974 && pixel_index <= 4976) || (pixel_index >= 4986 && pixel_index <= 4988) || (pixel_index >= 5000 && pixel_index <= 5006) || (pixel_index >= 5019 && pixel_index <= 5021) || (pixel_index >= 5031 && pixel_index <= 5043) || (pixel_index >= 5048 && pixel_index <= 5057) || (pixel_index >= 5070 && pixel_index <= 5072) || (pixel_index >= 5082 && pixel_index <= 5084) || (pixel_index >= 5096 && pixel_index <= 5102) || (pixel_index >= 5115 && pixel_index <= 5117) || (pixel_index >= 5127 && pixel_index <= 5139) || (pixel_index >= 5144 && pixel_index <= 5153) || (pixel_index >= 5166 && pixel_index <= 5168) || (pixel_index >= 5178 && pixel_index <= 5180) || (pixel_index >= 5192 && pixel_index <= 5198) || (pixel_index >= 5211 && pixel_index <= 5213) || (pixel_index >= 5223 && pixel_index <= 5235) || (pixel_index >= 5240 && pixel_index <= 5249) || (pixel_index >= 5262 && pixel_index <= 5264) || (pixel_index >= 5274 && pixel_index <= 5276) || (pixel_index >= 5295 && pixel_index <= 5297) || (pixel_index >= 5307 && pixel_index <= 5309) || (pixel_index >= 5319 && pixel_index <= 5321) || (pixel_index >= 5329 && pixel_index <= 5331) || (pixel_index >= 5336 && pixel_index <= 5338) || (pixel_index >= 5346 && pixel_index <= 5348) || (pixel_index >= 5358 && pixel_index <= 5360) || (pixel_index >= 5370 && pixel_index <= 5372) || (pixel_index >= 5381 && pixel_index <= 5383) || (pixel_index >= 5391 && pixel_index <= 5393) || (pixel_index >= 5403 && pixel_index <= 5405) || (pixel_index >= 5415 && pixel_index <= 5417) || (pixel_index >= 5425 && pixel_index <= 5427) || (pixel_index >= 5432 && pixel_index <= 5434) || (pixel_index >= 5442 && pixel_index <= 5444) || (pixel_index >= 5454 && pixel_index <= 5456) || (pixel_index >= 5477 && pixel_index <= 5479) || (pixel_index >= 5487 && pixel_index <= 5489) || (pixel_index >= 5499 && pixel_index <= 5501) || (pixel_index >= 5511 && pixel_index <= 5513) || (pixel_index >= 5521 && pixel_index <= 5523) || (pixel_index >= 5528 && pixel_index <= 5530) || (pixel_index >= 5538 && pixel_index <= 5540) || (pixel_index >= 5550 && pixel_index <= 5552) || (pixel_index >= 5573 && pixel_index <= 5575) || (pixel_index >= 5583 && pixel_index <= 5585) || (pixel_index >= 5595 && pixel_index <= 5597) || (pixel_index >= 5607 && pixel_index <= 5609) || (pixel_index >= 5617 && pixel_index <= 5619) || (pixel_index >= 5624 && pixel_index <= 5626) || (pixel_index >= 5634 && pixel_index <= 5636) || (pixel_index >= 5646 && pixel_index <= 5648) || (pixel_index >= 5669 && pixel_index <= 5671) || (pixel_index >= 5679 && pixel_index <= 5681) || (pixel_index >= 5691 && pixel_index <= 5693) || (pixel_index >= 5703 && pixel_index <= 5705) || (pixel_index >= 5713 && pixel_index <= 5715) || (pixel_index >= 5720 && pixel_index <= 5722) || (pixel_index >= 5730 && pixel_index <= 5732) || (pixel_index >= 5742 && pixel_index <= 5744) || (pixel_index >= 5768 && pixel_index <= 5774) || (pixel_index >= 5787 && pixel_index <= 5789) || (pixel_index >= 5799 && pixel_index <= 5801) || (pixel_index >= 5809 && pixel_index <= 5811) || (pixel_index >= 5816 && pixel_index <= 5818) || (pixel_index >= 5826 && pixel_index <= 5828) || (pixel_index >= 5838 && pixel_index <= 5840) || (pixel_index >= 5850 && pixel_index <= 5852) || (pixel_index >= 5864 && pixel_index <= 5870) || (pixel_index >= 5883 && pixel_index <= 5885) || (pixel_index >= 5895 && pixel_index <= 5897) || (pixel_index >= 5905 && pixel_index <= 5907) || (pixel_index >= 5912 && pixel_index <= 5914) || (pixel_index >= 5922 && pixel_index <= 5924) || (pixel_index >= 5934 && pixel_index <= 5936) || (pixel_index >= 5946 && pixel_index <= 5948) || (pixel_index >= 5960 && pixel_index <= 5966) || (pixel_index >= 5979 && pixel_index <= 5981) || (pixel_index >= 5991 && pixel_index <= 5993) || (pixel_index >= 6001 && pixel_index <= 6003) || (pixel_index >= 6008 && pixel_index <= 6010) || (pixel_index >= 6018 && pixel_index <= 6020) || (pixel_index >= 6030 && pixel_index <= 6032) || (pixel_index >= 6042 && pixel_index <= 6044)) begin
            oled_data = PINK_HEX;
        end else begin
            oled_data = BG_BLUE_HEX;
        end
    end
endmodule
