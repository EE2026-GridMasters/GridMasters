`timescale 1ns / 1ps

module display_winner(
    input clk,
    input [12:0] pixel_index,
    input [1:0] game_result,
    output [15:0] oled_data
    );

    wire [15:0] disp_winner_X, disp_winner_O, disp_draw;
    display_winner_X x (clk, pixel_index, disp_winner_X);
    display_winner_O o (clk, pixel_index, disp_winner_O);
    display_draw draw (clk, pixel_index, disp_draw);
    assign oled_data = (game_result == 2'b10) ? disp_winner_O :
        (game_result == 2'b01) ? disp_winner_X : disp_draw;
       
endmodule

module display_winner_X(
    input clk,
    input [12:0] pixel_index,
    output reg [15:0] oled_data
    );
    
    parameter PINK_HEX = 16'hF899;
    parameter BLUE_HEX = 16'h177F;
    parameter PURPLE_HEX = 16'h50DC;
    parameter BG_BLUE_HEX = 16'b0000000001000100;
    parameter WHITE_HEX = 16'hFFFF;
        
    wire anim_clk;
    custom_clock animclk (clk, 50_000_000, anim_clk);
    
    always @(clk) begin        
        if (anim_clk && ((pixel_index >= 635 && pixel_index <= 639) || (pixel_index >= 663 && pixel_index <= 667) || (pixel_index >= 731 && pixel_index <= 736) || (pixel_index >= 758 && pixel_index <= 763) || (pixel_index >= 827 && pixel_index <= 833) || (pixel_index >= 853 && pixel_index <= 859) || (pixel_index >= 923 && pixel_index <= 930) || (pixel_index >= 948 && pixel_index <= 955) || (pixel_index >= 1019 && pixel_index <= 1027) || (pixel_index >= 1043 && pixel_index <= 1051) || (pixel_index >= 1116 && pixel_index <= 1124) || (pixel_index >= 1138 && pixel_index <= 1146) || (pixel_index >= 1213 && pixel_index <= 1221) || (pixel_index >= 1233 && pixel_index <= 1241) || (pixel_index >= 1310 && pixel_index <= 1318) || (pixel_index >= 1328 && pixel_index <= 1336) || (pixel_index >= 1407 && pixel_index <= 1415) || (pixel_index >= 1423 && pixel_index <= 1431) || (pixel_index >= 1504 && pixel_index <= 1512) || (pixel_index >= 1518 && pixel_index <= 1526) || (pixel_index >= 1601 && pixel_index <= 1609) || (pixel_index >= 1613 && pixel_index <= 1621) || (pixel_index >= 1698 && pixel_index <= 1706) || (pixel_index >= 1708 && pixel_index <= 1716) || (pixel_index >= 1795 && pixel_index <= 1811) || (pixel_index >= 1892 && pixel_index <= 1906) || (pixel_index >= 1989 && pixel_index <= 2001) || (pixel_index >= 2086 && pixel_index <= 2096) || (pixel_index >= 2183 && pixel_index <= 2191) || (pixel_index >= 2226 && pixel_index <= 2228) || (pixel_index >= 2278 && pixel_index <= 2288) || (pixel_index >= 2322 && pixel_index <= 2324) || (pixel_index >= 2373 && pixel_index <= 2385) || (pixel_index >= 2418 && pixel_index <= 2420) || (pixel_index >= 2468 && pixel_index <= 2482) || (pixel_index >= 2514 && pixel_index <= 2516) || (pixel_index >= 2563 && pixel_index <= 2579) || (pixel_index >= 2610 && pixel_index <= 2612) || (pixel_index >= 2658 && pixel_index <= 2666) || (pixel_index >= 2668 && pixel_index <= 2676) || (pixel_index >= 2706 && pixel_index <= 2708) || (pixel_index >= 2753 && pixel_index <= 2761) || (pixel_index >= 2765 && pixel_index <= 2773) || (pixel_index >= 2798 && pixel_index <= 2808) || (pixel_index >= 2848 && pixel_index <= 2856) || (pixel_index >= 2862 && pixel_index <= 2870) || (pixel_index >= 2894 && pixel_index <= 2904) || (pixel_index >= 2943 && pixel_index <= 2951) || (pixel_index >= 2959 && pixel_index <= 2967) || (pixel_index >= 2990 && pixel_index <= 3000) || (pixel_index >= 3038 && pixel_index <= 3046) || (pixel_index >= 3056 && pixel_index <= 3064) || (pixel_index >= 3086 && pixel_index <= 3096) || (pixel_index >= 3133 && pixel_index <= 3141) || (pixel_index >= 3153 && pixel_index <= 3161) || (pixel_index >= 3175 && pixel_index <= 3199) || (pixel_index >= 3228 && pixel_index <= 3236) || (pixel_index >= 3250 && pixel_index <= 3258) || (pixel_index >= 3271 && pixel_index <= 3295) || (pixel_index >= 3324 && pixel_index <= 3331) || (pixel_index >= 3347 && pixel_index <= 3355) || (pixel_index >= 3367 && pixel_index <= 3391) || (pixel_index >= 3420 && pixel_index <= 3426) || (pixel_index >= 3444 && pixel_index <= 3451) || (pixel_index >= 3470 && pixel_index <= 3480) || (pixel_index >= 3516 && pixel_index <= 3521) || (pixel_index >= 3541 && pixel_index <= 3547) || (pixel_index >= 3566 && pixel_index <= 3576) || (pixel_index >= 3612 && pixel_index <= 3616) || (pixel_index >= 3638 && pixel_index <= 3643) || (pixel_index >= 3662 && pixel_index <= 3672) || (pixel_index >= 3735 && pixel_index <= 3739) || (pixel_index >= 3758 && pixel_index <= 3768) || (pixel_index >= 3858 && pixel_index <= 3860) || (pixel_index >= 3954 && pixel_index <= 3956) || (pixel_index >= 4050 && pixel_index <= 4052) || (pixel_index >= 4146 && pixel_index <= 4148) || (pixel_index >= 4242 && pixel_index <= 4244) || (pixel_index >= 4338 && pixel_index <= 4340))) begin
            oled_data <= BLUE_HEX;
        end else if (~anim_clk && ((pixel_index >= 635 && pixel_index <= 639) || (pixel_index >= 663 && pixel_index <= 667) || (pixel_index >= 731 && pixel_index <= 736) || (pixel_index >= 758 && pixel_index <= 763) || (pixel_index >= 827 && pixel_index <= 833) || (pixel_index >= 853 && pixel_index <= 859) || (pixel_index >= 923 && pixel_index <= 930) || (pixel_index >= 948 && pixel_index <= 955) || (pixel_index >= 1019 && pixel_index <= 1027) || (pixel_index >= 1043 && pixel_index <= 1051) || (pixel_index >= 1116 && pixel_index <= 1124) || (pixel_index >= 1138 && pixel_index <= 1146) || (pixel_index >= 1213 && pixel_index <= 1221) || (pixel_index >= 1233 && pixel_index <= 1241) || (pixel_index >= 1310 && pixel_index <= 1318) || (pixel_index >= 1328 && pixel_index <= 1336) || (pixel_index >= 1407 && pixel_index <= 1415) || (pixel_index >= 1423 && pixel_index <= 1431) || (pixel_index >= 1504 && pixel_index <= 1512) || (pixel_index >= 1518 && pixel_index <= 1526) || (pixel_index >= 1601 && pixel_index <= 1609) || (pixel_index >= 1613 && pixel_index <= 1621) || (pixel_index >= 1698 && pixel_index <= 1706) || (pixel_index >= 1708 && pixel_index <= 1716) || (pixel_index >= 1746 && pixel_index <= 1748) || (pixel_index >= 1795 && pixel_index <= 1811) || (pixel_index >= 1842 && pixel_index <= 1844) || (pixel_index >= 1892 && pixel_index <= 1906) || (pixel_index >= 1938 && pixel_index <= 1940) || (pixel_index >= 1989 && pixel_index <= 2001) || (pixel_index >= 2034 && pixel_index <= 2036) || (pixel_index >= 2086 && pixel_index <= 2096) || (pixel_index >= 2130 && pixel_index <= 2132) || (pixel_index >= 2183 && pixel_index <= 2191) || (pixel_index >= 2226 && pixel_index <= 2228) || (pixel_index >= 2278 && pixel_index <= 2288) || (pixel_index >= 2322 && pixel_index <= 2324) || (pixel_index >= 2373 && pixel_index <= 2385) || (pixel_index >= 2414 && pixel_index <= 2424) || (pixel_index >= 2468 && pixel_index <= 2482) || (pixel_index >= 2510 && pixel_index <= 2520) || (pixel_index >= 2563 && pixel_index <= 2579) || (pixel_index >= 2606 && pixel_index <= 2616) || (pixel_index >= 2658 && pixel_index <= 2666) || (pixel_index >= 2668 && pixel_index <= 2676) || (pixel_index >= 2702 && pixel_index <= 2712) || (pixel_index >= 2753 && pixel_index <= 2761) || (pixel_index >= 2765 && pixel_index <= 2773) || (pixel_index >= 2791 && pixel_index <= 2815) || (pixel_index >= 2848 && pixel_index <= 2856) || (pixel_index >= 2862 && pixel_index <= 2870) || (pixel_index >= 2887 && pixel_index <= 2911) || (pixel_index >= 2943 && pixel_index <= 2951) || (pixel_index >= 2959 && pixel_index <= 2967) || (pixel_index >= 2983 && pixel_index <= 3007) || (pixel_index >= 3038 && pixel_index <= 3046) || (pixel_index >= 3056 && pixel_index <= 3064) || (pixel_index >= 3086 && pixel_index <= 3096) || (pixel_index >= 3133 && pixel_index <= 3141) || (pixel_index >= 3153 && pixel_index <= 3161) || (pixel_index >= 3182 && pixel_index <= 3192) || (pixel_index >= 3228 && pixel_index <= 3236) || (pixel_index >= 3250 && pixel_index <= 3258) || (pixel_index >= 3278 && pixel_index <= 3288) || (pixel_index >= 3324 && pixel_index <= 3331) || (pixel_index >= 3347 && pixel_index <= 3355) || (pixel_index >= 3374 && pixel_index <= 3384) || (pixel_index >= 3420 && pixel_index <= 3426) || (pixel_index >= 3444 && pixel_index <= 3451) || (pixel_index >= 3474 && pixel_index <= 3476) || (pixel_index >= 3516 && pixel_index <= 3521) || (pixel_index >= 3541 && pixel_index <= 3547) || (pixel_index >= 3570 && pixel_index <= 3572) || (pixel_index >= 3612 && pixel_index <= 3616) || (pixel_index >= 3638 && pixel_index <= 3643) || (pixel_index >= 3666 && pixel_index <= 3668) || (pixel_index >= 3735 && pixel_index <= 3739) || (pixel_index >= 3762 && pixel_index <= 3764) || (pixel_index >= 3858 && pixel_index <= 3860) || (pixel_index >= 3954 && pixel_index <= 3956))) begin
            oled_data <= BLUE_HEX;
        end else if ((pixel_index >= 3969 && pixel_index <= 3971) || (pixel_index >= 3982 && pixel_index <= 3984) || (pixel_index >= 3989 && pixel_index <= 3991) || (pixel_index >= 3996 && pixel_index <= 3998) || (pixel_index >= 4009 && pixel_index <= 4011) || (pixel_index >= 4019 && pixel_index <= 4024) || (pixel_index >= 4065 && pixel_index <= 4067) || (pixel_index >= 4078 && pixel_index <= 4080) || (pixel_index >= 4085 && pixel_index <= 4087) || (pixel_index >= 4092 && pixel_index <= 4094) || (pixel_index >= 4105 && pixel_index <= 4107) || (pixel_index >= 4115 && pixel_index <= 4120) || (pixel_index >= 4161 && pixel_index <= 4163) || (pixel_index >= 4174 && pixel_index <= 4176) || (pixel_index >= 4181 && pixel_index <= 4183) || (pixel_index >= 4188 && pixel_index <= 4190) || (pixel_index >= 4201 && pixel_index <= 4203) || (pixel_index >= 4211 && pixel_index <= 4216) || (pixel_index >= 4257 && pixel_index <= 4259) || (pixel_index >= 4270 && pixel_index <= 4272) || (pixel_index >= 4277 && pixel_index <= 4279) || (pixel_index >= 4284 && pixel_index <= 4289) || (pixel_index >= 4297 && pixel_index <= 4299) || (pixel_index >= 4304 && pixel_index <= 4306) || (pixel_index >= 4313 && pixel_index <= 4315) || (pixel_index >= 4353 && pixel_index <= 4355) || (pixel_index >= 4366 && pixel_index <= 4368) || (pixel_index >= 4373 && pixel_index <= 4375) || (pixel_index >= 4380 && pixel_index <= 4385) || (pixel_index >= 4393 && pixel_index <= 4395) || (pixel_index >= 4400 && pixel_index <= 4402) || (pixel_index >= 4409 && pixel_index <= 4411) || (pixel_index >= 4449 && pixel_index <= 4451) || (pixel_index >= 4462 && pixel_index <= 4464) || (pixel_index >= 4469 && pixel_index <= 4471) || (pixel_index >= 4476 && pixel_index <= 4481) || (pixel_index >= 4489 && pixel_index <= 4491) || (pixel_index >= 4496 && pixel_index <= 4498) || (pixel_index >= 4505 && pixel_index <= 4507) || (pixel_index >= 4545 && pixel_index <= 4547) || (pixel_index >= 4552 && pixel_index <= 4554) || (pixel_index >= 4558 && pixel_index <= 4560) || (pixel_index >= 4565 && pixel_index <= 4567) || (pixel_index >= 4572 && pixel_index <= 4574) || (pixel_index >= 4578 && pixel_index <= 4580) || (pixel_index >= 4585 && pixel_index <= 4587) || (pixel_index >= 4592 && pixel_index <= 4594) || (pixel_index >= 4641 && pixel_index <= 4643) || (pixel_index >= 4648 && pixel_index <= 4650) || (pixel_index >= 4654 && pixel_index <= 4656) || (pixel_index >= 4661 && pixel_index <= 4663) || (pixel_index >= 4668 && pixel_index <= 4670) || (pixel_index >= 4674 && pixel_index <= 4676) || (pixel_index >= 4681 && pixel_index <= 4683) || (pixel_index >= 4691 && pixel_index <= 4696) || (pixel_index >= 4737 && pixel_index <= 4739) || (pixel_index >= 4744 && pixel_index <= 4746) || (pixel_index >= 4750 && pixel_index <= 4752) || (pixel_index >= 4757 && pixel_index <= 4759) || (pixel_index >= 4764 && pixel_index <= 4766) || (pixel_index >= 4770 && pixel_index <= 4772) || (pixel_index >= 4777 && pixel_index <= 4779) || (pixel_index >= 4787 && pixel_index <= 4792) || (pixel_index >= 4833 && pixel_index <= 4835) || (pixel_index >= 4840 && pixel_index <= 4842) || (pixel_index >= 4846 && pixel_index <= 4848) || (pixel_index >= 4853 && pixel_index <= 4855) || (pixel_index >= 4860 && pixel_index <= 4862) || (pixel_index >= 4869 && pixel_index <= 4875) || (pixel_index >= 4883 && pixel_index <= 4888) || (pixel_index >= 4929 && pixel_index <= 4931) || (pixel_index >= 4936 && pixel_index <= 4938) || (pixel_index >= 4942 && pixel_index <= 4944) || (pixel_index >= 4949 && pixel_index <= 4951) || (pixel_index >= 4956 && pixel_index <= 4958) || (pixel_index >= 4965 && pixel_index <= 4971) || (pixel_index >= 4985 && pixel_index <= 4987) || (pixel_index >= 5025 && pixel_index <= 5027) || (pixel_index >= 5032 && pixel_index <= 5034) || (pixel_index >= 5038 && pixel_index <= 5040) || (pixel_index >= 5045 && pixel_index <= 5047) || (pixel_index >= 5052 && pixel_index <= 5054) || (pixel_index >= 5061 && pixel_index <= 5067) || (pixel_index >= 5081 && pixel_index <= 5083) || (pixel_index >= 5121 && pixel_index <= 5127) || (pixel_index >= 5131 && pixel_index <= 5136) || (pixel_index >= 5141 && pixel_index <= 5143) || (pixel_index >= 5148 && pixel_index <= 5150) || (pixel_index >= 5161 && pixel_index <= 5163) || (pixel_index >= 5168 && pixel_index <= 5170) || (pixel_index >= 5177 && pixel_index <= 5179) || (pixel_index >= 5217 && pixel_index <= 5223) || (pixel_index >= 5227 && pixel_index <= 5232) || (pixel_index >= 5237 && pixel_index <= 5239) || (pixel_index >= 5244 && pixel_index <= 5246) || (pixel_index >= 5257 && pixel_index <= 5259) || (pixel_index >= 5264 && pixel_index <= 5266) || (pixel_index >= 5273 && pixel_index <= 5275) || (pixel_index >= 5313 && pixel_index <= 5319) || (pixel_index >= 5323 && pixel_index <= 5328) || (pixel_index >= 5333 && pixel_index <= 5335) || (pixel_index >= 5340 && pixel_index <= 5342) || (pixel_index >= 5353 && pixel_index <= 5355) || (pixel_index >= 5360 && pixel_index <= 5362) || (pixel_index >= 5369 && pixel_index <= 5371) || (pixel_index >= 5409 && pixel_index <= 5411) || (pixel_index >= 5422 && pixel_index <= 5424) || (pixel_index >= 5429 && pixel_index <= 5431) || (pixel_index >= 5436 && pixel_index <= 5438) || (pixel_index >= 5449 && pixel_index <= 5451) || (pixel_index >= 5459 && pixel_index <= 5464) || (pixel_index >= 5505 && pixel_index <= 5507) || (pixel_index >= 5518 && pixel_index <= 5520) || (pixel_index >= 5525 && pixel_index <= 5527) || (pixel_index >= 5532 && pixel_index <= 5534) || (pixel_index >= 5545 && pixel_index <= 5547) || (pixel_index >= 5555 && pixel_index <= 5560) || (pixel_index >= 5601 && pixel_index <= 5603) || (pixel_index >= 5614 && pixel_index <= 5616) || (pixel_index >= 5621 && pixel_index <= 5623) || (pixel_index >= 5628 && pixel_index <= 5630) || (pixel_index >= 5641 && pixel_index <= 5643) || (pixel_index >= 5651 && pixel_index <= 5656)) begin
            oled_data <= WHITE_HEX;
        end else begin
            oled_data <= BG_BLUE_HEX;
        end        
    end
endmodule

module display_winner_O(
    input clk,
    input [12:0] pixel_index,
    output reg [15:0] oled_data
    );
    parameter PINK_HEX = 16'hF899;
    parameter BLUE_HEX = 16'h177F;
    parameter PURPLE_HEX = 16'h50DC;
    parameter BG_BLUE_HEX = 16'h0006;
    parameter WHITE_HEX = 16'hFFFF;
    
    wire anim_clk;
    custom_clock animclk (clk, 50_000_000, anim_clk);
        
    always @(clk) begin
        if (anim_clk && ((pixel_index >= 646 && pixel_index <= 657) || (pixel_index >= 742 && pixel_index <= 753) || (pixel_index >= 833 && pixel_index <= 854) || (pixel_index >= 929 && pixel_index <= 950) || (pixel_index >= 1025 && pixel_index <= 1046) || (pixel_index >= 1119 && pixel_index <= 1128) || (pixel_index >= 1135 && pixel_index <= 1144) || (pixel_index >= 1215 && pixel_index <= 1224) || (pixel_index >= 1231 && pixel_index <= 1240) || (pixel_index >= 1311 && pixel_index <= 1315) || (pixel_index >= 1332 && pixel_index <= 1336) || (pixel_index >= 1407 && pixel_index <= 1411) || (pixel_index >= 1428 && pixel_index <= 1432) || (pixel_index >= 1503 && pixel_index <= 1507) || (pixel_index >= 1524 && pixel_index <= 1528) || (pixel_index >= 1596 && pixel_index <= 1603) || (pixel_index >= 1620 && pixel_index <= 1627) || (pixel_index >= 1692 && pixel_index <= 1699) || (pixel_index >= 1716 && pixel_index <= 1723) || (pixel_index >= 1788 && pixel_index <= 1792) || (pixel_index >= 1815 && pixel_index <= 1819) || (pixel_index >= 1884 && pixel_index <= 1888) || (pixel_index >= 1911 && pixel_index <= 1915) || (pixel_index >= 1980 && pixel_index <= 1984) || (pixel_index >= 2007 && pixel_index <= 2011) || (pixel_index >= 2076 && pixel_index <= 2080) || (pixel_index >= 2103 && pixel_index <= 2107) || (pixel_index >= 2130 && pixel_index <= 2132) || (pixel_index >= 2172 && pixel_index <= 2176) || (pixel_index >= 2199 && pixel_index <= 2203) || (pixel_index >= 2226 && pixel_index <= 2228) || (pixel_index >= 2268 && pixel_index <= 2272) || (pixel_index >= 2295 && pixel_index <= 2299) || (pixel_index >= 2322 && pixel_index <= 2324) || (pixel_index >= 2364 && pixel_index <= 2368) || (pixel_index >= 2391 && pixel_index <= 2395) || (pixel_index >= 2418 && pixel_index <= 2420) || (pixel_index >= 2460 && pixel_index <= 2467) || (pixel_index >= 2484 && pixel_index <= 2491) || (pixel_index >= 2514 && pixel_index <= 2516) || (pixel_index >= 2556 && pixel_index <= 2563) || (pixel_index >= 2580 && pixel_index <= 2587) || (pixel_index >= 2610 && pixel_index <= 2612) || (pixel_index >= 2652 && pixel_index <= 2659) || (pixel_index >= 2676 && pixel_index <= 2683) || (pixel_index >= 2706 && pixel_index <= 2708) || (pixel_index >= 2751 && pixel_index <= 2755) || (pixel_index >= 2772 && pixel_index <= 2776) || (pixel_index >= 2798 && pixel_index <= 2808) || (pixel_index >= 2847 && pixel_index <= 2851) || (pixel_index >= 2868 && pixel_index <= 2872) || (pixel_index >= 2894 && pixel_index <= 2904) || (pixel_index >= 2943 && pixel_index <= 2951) || (pixel_index >= 2960 && pixel_index <= 2968) || (pixel_index >= 2990 && pixel_index <= 3000) || (pixel_index >= 3039 && pixel_index <= 3047) || (pixel_index >= 3056 && pixel_index <= 3064) || (pixel_index >= 3086 && pixel_index <= 3096) || (pixel_index >= 3135 && pixel_index <= 3143) || (pixel_index >= 3152 && pixel_index <= 3160) || (pixel_index >= 3175 && pixel_index <= 3199) || (pixel_index >= 3233 && pixel_index <= 3254) || (pixel_index >= 3271 && pixel_index <= 3295) || (pixel_index >= 3329 && pixel_index <= 3350) || (pixel_index >= 3367 && pixel_index <= 3391) || (pixel_index >= 3429 && pixel_index <= 3442) || (pixel_index >= 3470 && pixel_index <= 3480) || (pixel_index >= 3525 && pixel_index <= 3538) || (pixel_index >= 3566 && pixel_index <= 3576) || (pixel_index >= 3621 && pixel_index <= 3634) || (pixel_index >= 3662 && pixel_index <= 3672) || (pixel_index >= 3758 && pixel_index <= 3768) || (pixel_index >= 3858 && pixel_index <= 3860) || (pixel_index >= 3954 && pixel_index <= 3956) || (pixel_index >= 4050 && pixel_index <= 4052) || (pixel_index >= 4146 && pixel_index <= 4148) || (pixel_index >= 4242 && pixel_index <= 4244) || (pixel_index >= 4338 && pixel_index <= 4340) || (pixel_index >= 4434 && pixel_index <= 4436))) begin
             oled_data <= PINK_HEX;
        end else if (~anim_clk && ((pixel_index >= 646 && pixel_index <= 657) || (pixel_index >= 742 && pixel_index <= 753) || (pixel_index >= 833 && pixel_index <= 854) || (pixel_index >= 929 && pixel_index <= 950) || (pixel_index >= 1025 && pixel_index <= 1046) || (pixel_index >= 1119 && pixel_index <= 1128) || (pixel_index >= 1135 && pixel_index <= 1144) || (pixel_index >= 1215 && pixel_index <= 1224) || (pixel_index >= 1231 && pixel_index <= 1240) || (pixel_index >= 1311 && pixel_index <= 1315) || (pixel_index >= 1332 && pixel_index <= 1336) || (pixel_index >= 1407 && pixel_index <= 1411) || (pixel_index >= 1428 && pixel_index <= 1432) || (pixel_index >= 1503 && pixel_index <= 1507) || (pixel_index >= 1524 && pixel_index <= 1528) || (pixel_index >= 1596 && pixel_index <= 1603) || (pixel_index >= 1620 && pixel_index <= 1627) || (pixel_index >= 1692 && pixel_index <= 1699) || (pixel_index >= 1716 && pixel_index <= 1723) || (pixel_index >= 1746 && pixel_index <= 1748) || (pixel_index >= 1788 && pixel_index <= 1792) || (pixel_index >= 1815 && pixel_index <= 1819) || (pixel_index >= 1842 && pixel_index <= 1844) || (pixel_index >= 1884 && pixel_index <= 1888) || (pixel_index >= 1911 && pixel_index <= 1915) || (pixel_index >= 1938 && pixel_index <= 1940) || (pixel_index >= 1980 && pixel_index <= 1984) || (pixel_index >= 2007 && pixel_index <= 2011) || (pixel_index >= 2034 && pixel_index <= 2036) || (pixel_index >= 2076 && pixel_index <= 2080) || (pixel_index >= 2103 && pixel_index <= 2107) || (pixel_index >= 2130 && pixel_index <= 2132) || (pixel_index >= 2172 && pixel_index <= 2176) || (pixel_index >= 2199 && pixel_index <= 2203) || (pixel_index >= 2226 && pixel_index <= 2228) || (pixel_index >= 2268 && pixel_index <= 2272) || (pixel_index >= 2295 && pixel_index <= 2299) || (pixel_index >= 2322 && pixel_index <= 2324) || (pixel_index >= 2364 && pixel_index <= 2368) || (pixel_index >= 2391 && pixel_index <= 2395) || (pixel_index >= 2414 && pixel_index <= 2424) || (pixel_index >= 2460 && pixel_index <= 2467) || (pixel_index >= 2484 && pixel_index <= 2491) || (pixel_index >= 2510 && pixel_index <= 2520) || (pixel_index >= 2556 && pixel_index <= 2563) || (pixel_index >= 2580 && pixel_index <= 2587) || (pixel_index >= 2606 && pixel_index <= 2616) || (pixel_index >= 2652 && pixel_index <= 2659) || (pixel_index >= 2676 && pixel_index <= 2683) || (pixel_index >= 2702 && pixel_index <= 2712) || (pixel_index >= 2751 && pixel_index <= 2755) || (pixel_index >= 2772 && pixel_index <= 2776) || (pixel_index >= 2791 && pixel_index <= 2815) || (pixel_index >= 2847 && pixel_index <= 2851) || (pixel_index >= 2868 && pixel_index <= 2872) || (pixel_index >= 2887 && pixel_index <= 2911) || (pixel_index >= 2943 && pixel_index <= 2951) || (pixel_index >= 2960 && pixel_index <= 2968) || (pixel_index >= 2983 && pixel_index <= 3007) || (pixel_index >= 3039 && pixel_index <= 3047) || (pixel_index >= 3056 && pixel_index <= 3064) || (pixel_index >= 3086 && pixel_index <= 3096) || (pixel_index >= 3135 && pixel_index <= 3143) || (pixel_index >= 3152 && pixel_index <= 3160) || (pixel_index >= 3182 && pixel_index <= 3192) || (pixel_index >= 3233 && pixel_index <= 3254) || (pixel_index >= 3278 && pixel_index <= 3288) || (pixel_index >= 3329 && pixel_index <= 3350) || (pixel_index >= 3374 && pixel_index <= 3384) || (pixel_index >= 3429 && pixel_index <= 3442) || (pixel_index >= 3474 && pixel_index <= 3476) || (pixel_index >= 3525 && pixel_index <= 3538) || (pixel_index >= 3570 && pixel_index <= 3572) || (pixel_index >= 3621 && pixel_index <= 3634) || (pixel_index >= 3666 && pixel_index <= 3668) || (pixel_index >= 3762 && pixel_index <= 3764) || (pixel_index >= 3858 && pixel_index <= 3860) || (pixel_index >= 3954 && pixel_index <= 3956))) begin
             oled_data <= PINK_HEX;
        end else if ((pixel_index >= 3969 && pixel_index <= 3971) || (pixel_index >= 3982 && pixel_index <= 3984) || (pixel_index >= 3989 && pixel_index <= 3991) || (pixel_index >= 3996 && pixel_index <= 3998) || (pixel_index >= 4009 && pixel_index <= 4011) || (pixel_index >= 4019 && pixel_index <= 4024) || (pixel_index >= 4065 && pixel_index <= 4067) || (pixel_index >= 4078 && pixel_index <= 4080) || (pixel_index >= 4085 && pixel_index <= 4087) || (pixel_index >= 4092 && pixel_index <= 4094) || (pixel_index >= 4105 && pixel_index <= 4107) || (pixel_index >= 4115 && pixel_index <= 4120) || (pixel_index >= 4161 && pixel_index <= 4163) || (pixel_index >= 4174 && pixel_index <= 4176) || (pixel_index >= 4181 && pixel_index <= 4183) || (pixel_index >= 4188 && pixel_index <= 4190) || (pixel_index >= 4201 && pixel_index <= 4203) || (pixel_index >= 4211 && pixel_index <= 4216) || (pixel_index >= 4257 && pixel_index <= 4259) || (pixel_index >= 4270 && pixel_index <= 4272) || (pixel_index >= 4277 && pixel_index <= 4279) || (pixel_index >= 4284 && pixel_index <= 4289) || (pixel_index >= 4297 && pixel_index <= 4299) || (pixel_index >= 4304 && pixel_index <= 4306) || (pixel_index >= 4313 && pixel_index <= 4315) || (pixel_index >= 4353 && pixel_index <= 4355) || (pixel_index >= 4366 && pixel_index <= 4368) || (pixel_index >= 4373 && pixel_index <= 4375) || (pixel_index >= 4380 && pixel_index <= 4385) || (pixel_index >= 4393 && pixel_index <= 4395) || (pixel_index >= 4400 && pixel_index <= 4402) || (pixel_index >= 4409 && pixel_index <= 4411) || (pixel_index >= 4449 && pixel_index <= 4451) || (pixel_index >= 4462 && pixel_index <= 4464) || (pixel_index >= 4469 && pixel_index <= 4471) || (pixel_index >= 4476 && pixel_index <= 4481) || (pixel_index >= 4489 && pixel_index <= 4491) || (pixel_index >= 4496 && pixel_index <= 4498) || (pixel_index >= 4505 && pixel_index <= 4507) || (pixel_index >= 4545 && pixel_index <= 4547) || (pixel_index >= 4552 && pixel_index <= 4554) || (pixel_index >= 4558 && pixel_index <= 4560) || (pixel_index >= 4565 && pixel_index <= 4567) || (pixel_index >= 4572 && pixel_index <= 4574) || (pixel_index >= 4578 && pixel_index <= 4580) || (pixel_index >= 4585 && pixel_index <= 4587) || (pixel_index >= 4592 && pixel_index <= 4594) || (pixel_index >= 4641 && pixel_index <= 4643) || (pixel_index >= 4648 && pixel_index <= 4650) || (pixel_index >= 4654 && pixel_index <= 4656) || (pixel_index >= 4661 && pixel_index <= 4663) || (pixel_index >= 4668 && pixel_index <= 4670) || (pixel_index >= 4674 && pixel_index <= 4676) || (pixel_index >= 4681 && pixel_index <= 4683) || (pixel_index >= 4691 && pixel_index <= 4696) || (pixel_index >= 4737 && pixel_index <= 4739) || (pixel_index >= 4744 && pixel_index <= 4746) || (pixel_index >= 4750 && pixel_index <= 4752) || (pixel_index >= 4757 && pixel_index <= 4759) || (pixel_index >= 4764 && pixel_index <= 4766) || (pixel_index >= 4770 && pixel_index <= 4772) || (pixel_index >= 4777 && pixel_index <= 4779) || (pixel_index >= 4787 && pixel_index <= 4792) || (pixel_index >= 4833 && pixel_index <= 4835) || (pixel_index >= 4840 && pixel_index <= 4842) || (pixel_index >= 4846 && pixel_index <= 4848) || (pixel_index >= 4853 && pixel_index <= 4855) || (pixel_index >= 4860 && pixel_index <= 4862) || (pixel_index >= 4869 && pixel_index <= 4875) || (pixel_index >= 4883 && pixel_index <= 4888) || (pixel_index >= 4929 && pixel_index <= 4931) || (pixel_index >= 4936 && pixel_index <= 4938) || (pixel_index >= 4942 && pixel_index <= 4944) || (pixel_index >= 4949 && pixel_index <= 4951) || (pixel_index >= 4956 && pixel_index <= 4958) || (pixel_index >= 4965 && pixel_index <= 4971) || (pixel_index >= 4985 && pixel_index <= 4987) || (pixel_index >= 5025 && pixel_index <= 5027) || (pixel_index >= 5032 && pixel_index <= 5034) || (pixel_index >= 5038 && pixel_index <= 5040) || (pixel_index >= 5045 && pixel_index <= 5047) || (pixel_index >= 5052 && pixel_index <= 5054) || (pixel_index >= 5061 && pixel_index <= 5067) || (pixel_index >= 5081 && pixel_index <= 5083) || (pixel_index >= 5121 && pixel_index <= 5127) || (pixel_index >= 5131 && pixel_index <= 5136) || (pixel_index >= 5141 && pixel_index <= 5143) || (pixel_index >= 5148 && pixel_index <= 5150) || (pixel_index >= 5161 && pixel_index <= 5163) || (pixel_index >= 5168 && pixel_index <= 5170) || (pixel_index >= 5177 && pixel_index <= 5179) || (pixel_index >= 5217 && pixel_index <= 5223) || (pixel_index >= 5227 && pixel_index <= 5232) || (pixel_index >= 5237 && pixel_index <= 5239) || (pixel_index >= 5244 && pixel_index <= 5246) || (pixel_index >= 5257 && pixel_index <= 5259) || (pixel_index >= 5264 && pixel_index <= 5266) || (pixel_index >= 5273 && pixel_index <= 5275) || (pixel_index >= 5313 && pixel_index <= 5319) || (pixel_index >= 5323 && pixel_index <= 5328) || (pixel_index >= 5333 && pixel_index <= 5335) || (pixel_index >= 5340 && pixel_index <= 5342) || (pixel_index >= 5353 && pixel_index <= 5355) || (pixel_index >= 5360 && pixel_index <= 5362) || (pixel_index >= 5369 && pixel_index <= 5371) || (pixel_index >= 5409 && pixel_index <= 5411) || (pixel_index >= 5422 && pixel_index <= 5424) || (pixel_index >= 5429 && pixel_index <= 5431) || (pixel_index >= 5436 && pixel_index <= 5438) || (pixel_index >= 5449 && pixel_index <= 5451) || (pixel_index >= 5459 && pixel_index <= 5464) || (pixel_index >= 5505 && pixel_index <= 5507) || (pixel_index >= 5518 && pixel_index <= 5520) || (pixel_index >= 5525 && pixel_index <= 5527) || (pixel_index >= 5532 && pixel_index <= 5534) || (pixel_index >= 5545 && pixel_index <= 5547) || (pixel_index >= 5555 && pixel_index <= 5560) || (pixel_index >= 5601 && pixel_index <= 5603) || (pixel_index >= 5614 && pixel_index <= 5616) || (pixel_index >= 5621 && pixel_index <= 5623) || (pixel_index >= 5628 && pixel_index <= 5630) || (pixel_index >= 5641 && pixel_index <= 5643) || (pixel_index >= 5651 && pixel_index <= 5656)) begin
            oled_data <= WHITE_HEX;
        end else begin
            oled_data <= BG_BLUE_HEX;
        end
    end
endmodule

module display_draw(
    input clk,
    input [12:0] pixel_index,
    output reg [15:0] oled_data
    );
    
    parameter PINK_HEX = 16'hF899;
    parameter BLUE_HEX = 16'h177F;
    parameter BG_BLUE_HEX = 16'h0006;
    parameter WHITE_HEX = 16'hFFFF;
    
    always @(*) begin
        if ((pixel_index >= 641 && pixel_index <= 648) || (pixel_index >= 734 && pixel_index <= 746) || (pixel_index >= 828 && pixel_index <= 844) || (pixel_index >= 922 && pixel_index <= 927) || (pixel_index >= 937 && pixel_index <= 942) || (pixel_index >= 1017 && pixel_index <= 1021) || (pixel_index >= 1035 && pixel_index <= 1039) || (pixel_index >= 1112 && pixel_index <= 1115) || (pixel_index >= 1132 && pixel_index <= 1136) || (pixel_index >= 1207 && pixel_index <= 1210) || (pixel_index >= 1230 && pixel_index <= 1233) || (pixel_index >= 1302 && pixel_index <= 1305) || (pixel_index >= 1327 && pixel_index <= 1330) || (pixel_index >= 1398 && pixel_index <= 1401) || (pixel_index >= 1424 && pixel_index <= 1426) || (pixel_index >= 1493 && pixel_index <= 1496) || (pixel_index >= 1520 && pixel_index <= 1523) || (pixel_index >= 1589 && pixel_index <= 1592) || (pixel_index >= 1617 && pixel_index <= 1619) || (pixel_index >= 1685 && pixel_index <= 1687) || (pixel_index >= 1713 && pixel_index <= 1715) || (pixel_index >= 1780 && pixel_index <= 1783) || (pixel_index >= 1810 && pixel_index <= 1812) || (pixel_index >= 1876 && pixel_index <= 1878) || (pixel_index >= 1906 && pixel_index <= 1908) || (pixel_index >= 1972 && pixel_index <= 1974) || (pixel_index >= 2002 && pixel_index <= 2004) || (pixel_index >= 2068 && pixel_index <= 2070) || (pixel_index >= 2098 && pixel_index <= 2100) || (pixel_index >= 2164 && pixel_index <= 2166) || (pixel_index >= 2194 && pixel_index <= 2196) || (pixel_index >= 2260 && pixel_index <= 2262) || (pixel_index >= 2290 && pixel_index <= 2292) || (pixel_index >= 2356 && pixel_index <= 2359) || (pixel_index >= 2385 && pixel_index <= 2388) || (pixel_index >= 2453 && pixel_index <= 2455) || (pixel_index >= 2481 && pixel_index <= 2483) || (pixel_index >= 2549 && pixel_index <= 2552) || (pixel_index >= 2577 && pixel_index <= 2579) || (pixel_index >= 2645 && pixel_index <= 2648) || (pixel_index >= 2672 && pixel_index <= 2675) || (pixel_index >= 2742 && pixel_index <= 2745) || (pixel_index >= 2768 && pixel_index <= 2770) || (pixel_index >= 2838 && pixel_index <= 2841) || (pixel_index >= 2863 && pixel_index <= 2866) || (pixel_index >= 2935 && pixel_index <= 2938) || (pixel_index >= 2957 && pixel_index <= 2961) || (pixel_index >= 3032 && pixel_index <= 3036) || (pixel_index >= 3052 && pixel_index <= 3056) || (pixel_index >= 3129 && pixel_index <= 3134) || (pixel_index >= 3146 && pixel_index <= 3151) || (pixel_index >= 3226 && pixel_index <= 3232) || (pixel_index >= 3240 && pixel_index <= 3246) || (pixel_index >= 3324 && pixel_index <= 3340) || (pixel_index >= 3422 && pixel_index <= 3434) || (pixel_index >= 3521 && pixel_index <= 3527)) begin
            oled_data = PINK_HEX;
        end else if ((pixel_index >= 684 && pixel_index <= 688) || (pixel_index >= 710 && pixel_index <= 713) || (pixel_index >= 780 && pixel_index <= 785) || (pixel_index >= 805 && pixel_index <= 809) || (pixel_index >= 876 && pixel_index <= 882) || (pixel_index >= 900 && pixel_index <= 905) || (pixel_index >= 972 && pixel_index <= 979) || (pixel_index >= 995 && pixel_index <= 1001) || (pixel_index >= 1069 && pixel_index <= 1076) || (pixel_index >= 1090 && pixel_index <= 1096) || (pixel_index >= 1166 && pixel_index <= 1173) || (pixel_index >= 1185 && pixel_index <= 1191) || (pixel_index >= 1263 && pixel_index <= 1270) || (pixel_index >= 1280 && pixel_index <= 1286) || (pixel_index >= 1360 && pixel_index <= 1367) || (pixel_index >= 1375 && pixel_index <= 1381) || (pixel_index >= 1457 && pixel_index <= 1464) || (pixel_index >= 1470 && pixel_index <= 1476) || (pixel_index >= 1554 && pixel_index <= 1561) || (pixel_index >= 1565 && pixel_index <= 1571) || (pixel_index >= 1651 && pixel_index <= 1658) || (pixel_index >= 1660 && pixel_index <= 1666) || (pixel_index >= 1748 && pixel_index <= 1761) || (pixel_index >= 1845 && pixel_index <= 1856) || (pixel_index >= 1942 && pixel_index <= 1951) || (pixel_index >= 2039 && pixel_index <= 2046) || (pixel_index >= 2135 && pixel_index <= 2142) || (pixel_index >= 2230 && pixel_index <= 2239) || (pixel_index >= 2325 && pixel_index <= 2336) || (pixel_index >= 2420 && pixel_index <= 2433) || (pixel_index >= 2515 && pixel_index <= 2521) || (pixel_index >= 2524 && pixel_index <= 2530) || (pixel_index >= 2610 && pixel_index <= 2616) || (pixel_index >= 2621 && pixel_index <= 2627) || (pixel_index >= 2705 && pixel_index <= 2711) || (pixel_index >= 2718 && pixel_index <= 2724) || (pixel_index >= 2800 && pixel_index <= 2806) || (pixel_index >= 2815 && pixel_index <= 2821) || (pixel_index >= 2895 && pixel_index <= 2901) || (pixel_index >= 2912 && pixel_index <= 2918) || (pixel_index >= 2990 && pixel_index <= 2996) || (pixel_index >= 3009 && pixel_index <= 3015) || (pixel_index >= 3085 && pixel_index <= 3091) || (pixel_index >= 3106 && pixel_index <= 3112) || (pixel_index >= 3180 && pixel_index <= 3186) || (pixel_index >= 3203 && pixel_index <= 3209) || (pixel_index >= 3276 && pixel_index <= 3281) || (pixel_index >= 3300 && pixel_index <= 3305) || (pixel_index >= 3372 && pixel_index <= 3376) || (pixel_index >= 3397 && pixel_index <= 3401) || (pixel_index >= 3468 && pixel_index <= 3471) || (pixel_index >= 3494 && pixel_index <= 3497)) begin
            oled_data = BLUE_HEX;
        end else if ((pixel_index >= 3856 && pixel_index <= 3864) || (pixel_index >= 3872 && pixel_index <= 3880) || (pixel_index >= 3891 && pixel_index <= 3897) || (pixel_index >= 3905 && pixel_index <= 3907) || (pixel_index >= 3918 && pixel_index <= 3920) || (pixel_index >= 3952 && pixel_index <= 3960) || (pixel_index >= 3968 && pixel_index <= 3976) || (pixel_index >= 3987 && pixel_index <= 3993) || (pixel_index >= 4001 && pixel_index <= 4003) || (pixel_index >= 4014 && pixel_index <= 4016) || (pixel_index >= 4048 && pixel_index <= 4056) || (pixel_index >= 4064 && pixel_index <= 4072) || (pixel_index >= 4083 && pixel_index <= 4089) || (pixel_index >= 4097 && pixel_index <= 4099) || (pixel_index >= 4110 && pixel_index <= 4112) || (pixel_index >= 4144 && pixel_index <= 4146) || (pixel_index >= 4153 && pixel_index <= 4155) || (pixel_index >= 4160 && pixel_index <= 4162) || (pixel_index >= 4169 && pixel_index <= 4171) || (pixel_index >= 4176 && pixel_index <= 4178) || (pixel_index >= 4186 && pixel_index <= 4188) || (pixel_index >= 4193 && pixel_index <= 4195) || (pixel_index >= 4206 && pixel_index <= 4208) || (pixel_index >= 4240 && pixel_index <= 4242) || (pixel_index >= 4249 && pixel_index <= 4251) || (pixel_index >= 4256 && pixel_index <= 4258) || (pixel_index >= 4265 && pixel_index <= 4267) || (pixel_index >= 4272 && pixel_index <= 4274) || (pixel_index >= 4282 && pixel_index <= 4284) || (pixel_index >= 4289 && pixel_index <= 4291) || (pixel_index >= 4302 && pixel_index <= 4304) || (pixel_index >= 4336 && pixel_index <= 4338) || (pixel_index >= 4345 && pixel_index <= 4347) || (pixel_index >= 4352 && pixel_index <= 4354) || (pixel_index >= 4361 && pixel_index <= 4363) || (pixel_index >= 4368 && pixel_index <= 4370) || (pixel_index >= 4378 && pixel_index <= 4380) || (pixel_index >= 4385 && pixel_index <= 4387) || (pixel_index >= 4398 && pixel_index <= 4400) || (pixel_index >= 4432 && pixel_index <= 4434) || (pixel_index >= 4441 && pixel_index <= 4443) || (pixel_index >= 4448 && pixel_index <= 4450) || (pixel_index >= 4457 && pixel_index <= 4459) || (pixel_index >= 4464 && pixel_index <= 4466) || (pixel_index >= 4474 && pixel_index <= 4476) || (pixel_index >= 4481 && pixel_index <= 4483) || (pixel_index >= 4487 && pixel_index <= 4489) || (pixel_index >= 4494 && pixel_index <= 4496) || (pixel_index >= 4528 && pixel_index <= 4530) || (pixel_index >= 4537 && pixel_index <= 4539) || (pixel_index >= 4544 && pixel_index <= 4546) || (pixel_index >= 4553 && pixel_index <= 4555) || (pixel_index >= 4560 && pixel_index <= 4562) || (pixel_index >= 4570 && pixel_index <= 4572) || (pixel_index >= 4577 && pixel_index <= 4579) || (pixel_index >= 4583 && pixel_index <= 4585) || (pixel_index >= 4590 && pixel_index <= 4592) || (pixel_index >= 4624 && pixel_index <= 4626) || (pixel_index >= 4633 && pixel_index <= 4635) || (pixel_index >= 4640 && pixel_index <= 4648) || (pixel_index >= 4656 && pixel_index <= 4668) || (pixel_index >= 4673 && pixel_index <= 4675) || (pixel_index >= 4679 && pixel_index <= 4681) || (pixel_index >= 4686 && pixel_index <= 4688) || (pixel_index >= 4720 && pixel_index <= 4722) || (pixel_index >= 4729 && pixel_index <= 4731) || (pixel_index >= 4736 && pixel_index <= 4744) || (pixel_index >= 4752 && pixel_index <= 4764) || (pixel_index >= 4769 && pixel_index <= 4771) || (pixel_index >= 4775 && pixel_index <= 4777) || (pixel_index >= 4782 && pixel_index <= 4784) || (pixel_index >= 4816 && pixel_index <= 4818) || (pixel_index >= 4825 && pixel_index <= 4827) || (pixel_index >= 4832 && pixel_index <= 4840) || (pixel_index >= 4848 && pixel_index <= 4860) || (pixel_index >= 4865 && pixel_index <= 4867) || (pixel_index >= 4871 && pixel_index <= 4873) || (pixel_index >= 4878 && pixel_index <= 4880) || (pixel_index >= 4912 && pixel_index <= 4914) || (pixel_index >= 4921 && pixel_index <= 4923) || (pixel_index >= 4928 && pixel_index <= 4930) || (pixel_index >= 4937 && pixel_index <= 4939) || (pixel_index >= 4944 && pixel_index <= 4946) || (pixel_index >= 4954 && pixel_index <= 4956) || (pixel_index >= 4961 && pixel_index <= 4963) || (pixel_index >= 4967 && pixel_index <= 4969) || (pixel_index >= 4974 && pixel_index <= 4976) || (pixel_index >= 5008 && pixel_index <= 5010) || (pixel_index >= 5017 && pixel_index <= 5019) || (pixel_index >= 5024 && pixel_index <= 5026) || (pixel_index >= 5033 && pixel_index <= 5035) || (pixel_index >= 5040 && pixel_index <= 5042) || (pixel_index >= 5050 && pixel_index <= 5052) || (pixel_index >= 5057 && pixel_index <= 5062) || (pixel_index >= 5066 && pixel_index <= 5072) || (pixel_index >= 5104 && pixel_index <= 5106) || (pixel_index >= 5113 && pixel_index <= 5115) || (pixel_index >= 5120 && pixel_index <= 5122) || (pixel_index >= 5129 && pixel_index <= 5131) || (pixel_index >= 5136 && pixel_index <= 5138) || (pixel_index >= 5146 && pixel_index <= 5148) || (pixel_index >= 5153 && pixel_index <= 5158) || (pixel_index >= 5162 && pixel_index <= 5168) || (pixel_index >= 5200 && pixel_index <= 5202) || (pixel_index >= 5209 && pixel_index <= 5211) || (pixel_index >= 5216 && pixel_index <= 5218) || (pixel_index >= 5225 && pixel_index <= 5227) || (pixel_index >= 5232 && pixel_index <= 5234) || (pixel_index >= 5242 && pixel_index <= 5244) || (pixel_index >= 5249 && pixel_index <= 5254) || (pixel_index >= 5258 && pixel_index <= 5264) || (pixel_index >= 5296 && pixel_index <= 5298) || (pixel_index >= 5305 && pixel_index <= 5307) || (pixel_index >= 5312 && pixel_index <= 5314) || (pixel_index >= 5321 && pixel_index <= 5323) || (pixel_index >= 5328 && pixel_index <= 5330) || (pixel_index >= 5338 && pixel_index <= 5340) || (pixel_index >= 5345 && pixel_index <= 5347) || (pixel_index >= 5358 && pixel_index <= 5360) || (pixel_index >= 5392 && pixel_index <= 5400) || (pixel_index >= 5408 && pixel_index <= 5410) || (pixel_index >= 5417 && pixel_index <= 5419) || (pixel_index >= 5424 && pixel_index <= 5426) || (pixel_index >= 5434 && pixel_index <= 5436) || (pixel_index >= 5441 && pixel_index <= 5443) || (pixel_index >= 5454 && pixel_index <= 5456) || (pixel_index >= 5488 && pixel_index <= 5496) || (pixel_index >= 5504 && pixel_index <= 5506) || (pixel_index >= 5513 && pixel_index <= 5515) || (pixel_index >= 5520 && pixel_index <= 5522) || (pixel_index >= 5530 && pixel_index <= 5532) || (pixel_index >= 5537 && pixel_index <= 5539) || (pixel_index >= 5550 && pixel_index <= 5552) || (pixel_index >= 5584 && pixel_index <= 5592) || (pixel_index >= 5600 && pixel_index <= 5602) || (pixel_index >= 5609 && pixel_index <= 5611) || (pixel_index >= 5616 && pixel_index <= 5618) || (pixel_index >= 5626 && pixel_index <= 5628) || (pixel_index >= 5633 && pixel_index <= 5635) || (pixel_index >= 5646 && pixel_index <= 5648)) begin
            oled_data = WHITE_HEX;
        end else begin
            oled_data = BG_BLUE_HEX;
        end
    end
    
endmodule