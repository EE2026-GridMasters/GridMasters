`timescale 1ns / 1ps

module combase_data(input [12:0] pixel_index, output reg [15:0] oled_data);
   
    always @ (*) begin
        if (((pixel_index >= 194) && (pixel_index <= 285)) || ((pixel_index >= 290) && (pixel_index <= 381)) || ((pixel_index >= 386) && (pixel_index <= 387)) || ((pixel_index >= 476) && (pixel_index <= 477)) || ((pixel_index >= 482) && (pixel_index <= 483)) || ((pixel_index >= 572) && (pixel_index <= 573)) || ((pixel_index >= 578) && (pixel_index <= 579)) || ((pixel_index >= 600) && (pixel_index <= 601)) || ((pixel_index >= 608) && (pixel_index <= 609)) || ((pixel_index >= 614) && (pixel_index <= 619)) || ((pixel_index >= 636) && (pixel_index <= 639)) || ((pixel_index >= 644) && (pixel_index <= 649)) || ((pixel_index >= 668) && (pixel_index <= 669)) || ((pixel_index >= 674) && (pixel_index <= 675)) || ((pixel_index >= 696) && (pixel_index <= 697)) || ((pixel_index >= 704) && (pixel_index <= 705)) || ((pixel_index >= 710) && (pixel_index <= 715)) || ((pixel_index >= 732) && (pixel_index <= 735)) || ((pixel_index >= 740) && (pixel_index <= 745)) || ((pixel_index >= 764) && (pixel_index <= 765)) || ((pixel_index >= 770) && (pixel_index <= 771)) || ((pixel_index >= 792) && (pixel_index <= 793)) || ((pixel_index >= 800) && (pixel_index <= 801)) || ((pixel_index >= 804) && (pixel_index <= 805)) || ((pixel_index >= 826) && (pixel_index <= 827)) || ((pixel_index >= 832) && (pixel_index <= 833)) || ((pixel_index >= 838) && (pixel_index <= 839)) || ((pixel_index >= 860) && (pixel_index <= 861)) || ((pixel_index >= 866) && (pixel_index <= 867)) || ((pixel_index >= 888) && (pixel_index <= 889)) || ((pixel_index >= 896) && (pixel_index <= 897)) || ((pixel_index >= 900) && (pixel_index <= 901)) || ((pixel_index >= 922) && (pixel_index <= 923)) || ((pixel_index >= 928) && (pixel_index <= 929)) || ((pixel_index >= 934) && (pixel_index <= 935)) || ((pixel_index >= 956) && (pixel_index <= 957)) || ((pixel_index >= 962) && (pixel_index <= 963)) || ((pixel_index >= 986) && (pixel_index <= 987)) || ((pixel_index >= 990) && (pixel_index <= 991)) || ((pixel_index >= 998) && (pixel_index <= 1001)) || ((pixel_index >= 1018) && (pixel_index <= 1025)) || ((pixel_index >= 1030) && (pixel_index <= 1031)) || ((pixel_index >= 1052) && (pixel_index <= 1053)) || ((pixel_index >= 1058) && (pixel_index <= 1059)) || ((pixel_index >= 1082) && (pixel_index <= 1083)) || ((pixel_index >= 1086) && (pixel_index <= 1087)) || ((pixel_index >= 1094) && (pixel_index <= 1097)) || ((pixel_index >= 1114) && (pixel_index <= 1121)) || ((pixel_index >= 1126) && (pixel_index <= 1127)) || ((pixel_index >= 1148) && (pixel_index <= 1149)) || ((pixel_index >= 1154) && (pixel_index <= 1155)) || ((pixel_index >= 1178) && (pixel_index <= 1179)) || ((pixel_index >= 1182) && (pixel_index <= 1183)) || ((pixel_index >= 1194) && (pixel_index <= 1195)) || ((pixel_index >= 1210) && (pixel_index <= 1211)) || ((pixel_index >= 1216) && (pixel_index <= 1217)) || ((pixel_index >= 1222) && (pixel_index <= 1223)) || ((pixel_index >= 1244) && (pixel_index <= 1245)) || ((pixel_index >= 1250) && (pixel_index <= 1251)) || ((pixel_index >= 1274) && (pixel_index <= 1275)) || ((pixel_index >= 1278) && (pixel_index <= 1279)) || ((pixel_index >= 1290) && (pixel_index <= 1291)) || ((pixel_index >= 1306) && (pixel_index <= 1307)) || ((pixel_index >= 1312) && (pixel_index <= 1313)) || ((pixel_index >= 1318) && (pixel_index <= 1319)) || ((pixel_index >= 1340) && (pixel_index <= 1341)) || ((pixel_index >= 1346) && (pixel_index <= 1347)) || ((pixel_index >= 1372) && (pixel_index <= 1373)) || ((pixel_index >= 1380) && (pixel_index <= 1385)) || ((pixel_index >= 1392) && (pixel_index <= 1393)) || ((pixel_index >= 1402) && (pixel_index <= 1403)) || ((pixel_index >= 1408) && (pixel_index <= 1409)) || ((pixel_index >= 1412) && (pixel_index <= 1417)) || ((pixel_index >= 1436) && (pixel_index <= 1437)) || ((pixel_index >= 1442) && (pixel_index <= 1443)) || ((pixel_index >= 1468) && (pixel_index <= 1469)) || ((pixel_index >= 1476) && (pixel_index <= 1481)) || ((pixel_index >= 1488) && (pixel_index <= 1489)) || ((pixel_index >= 1498) && (pixel_index <= 1499)) || ((pixel_index >= 1504) && (pixel_index <= 1505)) || ((pixel_index >= 1508) && (pixel_index <= 1513)) || ((pixel_index >= 1532) && (pixel_index <= 1533)) || ((pixel_index >= 1538) && (pixel_index <= 1539)) || ((pixel_index >= 1628) && (pixel_index <= 1629)) || ((pixel_index >= 1634) && (pixel_index <= 1635)) || ((pixel_index >= 1724) && (pixel_index <= 1725)) || ((pixel_index >= 1730) && (pixel_index <= 1821)) || ((pixel_index >= 1826) && (pixel_index <= 1917)) || ((pixel_index >= 2232) && (pixel_index <= 2233)) || ((pixel_index >= 2242) && (pixel_index <= 2249)) || ((pixel_index >= 2252) && (pixel_index <= 2253)) || ((pixel_index >= 2260) && (pixel_index <= 2261)) || ((pixel_index >= 2264) && (pixel_index <= 2271)) || ((pixel_index >= 2274) && (pixel_index <= 2275)) || ((pixel_index >= 2328) && (pixel_index <= 2329)) || ((pixel_index >= 2338) && (pixel_index <= 2345)) || ((pixel_index >= 2348) && (pixel_index <= 2349)) || ((pixel_index >= 2356) && (pixel_index <= 2357)) || ((pixel_index >= 2360) && (pixel_index <= 2367)) || ((pixel_index >= 2370) && (pixel_index <= 2371)) || ((pixel_index >= 2424) && (pixel_index <= 2425)) || ((pixel_index >= 2434) && (pixel_index <= 2435)) || ((pixel_index >= 2444) && (pixel_index <= 2445)) || ((pixel_index >= 2452) && (pixel_index <= 2453)) || ((pixel_index >= 2456) && (pixel_index <= 2457)) || ((pixel_index >= 2466) && (pixel_index <= 2467)) || ((pixel_index >= 2520) && (pixel_index <= 2521)) || ((pixel_index >= 2530) && (pixel_index <= 2531)) || ((pixel_index >= 2540) && (pixel_index <= 2541)) || ((pixel_index >= 2548) && (pixel_index <= 2549)) || ((pixel_index >= 2552) && (pixel_index <= 2553)) || ((pixel_index >= 2562) && (pixel_index <= 2563)) || ((pixel_index >= 2616) && (pixel_index <= 2617)) || ((pixel_index >= 2626) && (pixel_index <= 2631)) || ((pixel_index >= 2638) && (pixel_index <= 2639)) || ((pixel_index >= 2642) && (pixel_index <= 2643)) || ((pixel_index >= 2648) && (pixel_index <= 2653)) || ((pixel_index >= 2658) && (pixel_index <= 2659)) || ((pixel_index >= 2712) && (pixel_index <= 2713)) || ((pixel_index >= 2722) && (pixel_index <= 2727)) || ((pixel_index >= 2734) && (pixel_index <= 2735)) || ((pixel_index >= 2738) && (pixel_index <= 2739)) || ((pixel_index >= 2744) && (pixel_index <= 2749)) || ((pixel_index >= 2754) && (pixel_index <= 2755)) || ((pixel_index >= 2808) && (pixel_index <= 2809)) || ((pixel_index >= 2818) && (pixel_index <= 2819)) || ((pixel_index >= 2830) && (pixel_index <= 2831)) || ((pixel_index >= 2834) && (pixel_index <= 2835)) || ((pixel_index >= 2840) && (pixel_index <= 2841)) || ((pixel_index >= 2850) && (pixel_index <= 2851)) || ((pixel_index >= 2904) && (pixel_index <= 2905)) || ((pixel_index >= 2914) && (pixel_index <= 2915)) || ((pixel_index >= 2926) && (pixel_index <= 2927)) || ((pixel_index >= 2930) && (pixel_index <= 2931)) || ((pixel_index >= 2936) && (pixel_index <= 2937)) || ((pixel_index >= 2946) && (pixel_index <= 2947)) || ((pixel_index >= 3000) && (pixel_index <= 3007)) || ((pixel_index >= 3010) && (pixel_index <= 3017)) || ((pixel_index >= 3024) && (pixel_index <= 3025)) || ((pixel_index >= 3032) && (pixel_index <= 3039)) || ((pixel_index >= 3042) && (pixel_index <= 3049)) || ((pixel_index >= 3096) && (pixel_index <= 3103)) || ((pixel_index >= 3106) && (pixel_index <= 3113)) || ((pixel_index >= 3120) && (pixel_index <= 3121)) || ((pixel_index >= 3128) && (pixel_index <= 3135)) || (pixel_index >= 3138) && (pixel_index <= 3145)) oled_data = 16'b1111111111111111;
        else if (pixel_index >= 3264) oled_data = 0;
        else oled_data = 16'b0000000001000100;
    end

endmodule

module comlvl_data(input [1:0] sw, input [12:0] pixel_index, output reg [15:0] oled_data);
    wire [6:0] x = pixel_index % 96;
    wire [6:0] y = pixel_index / 96;
   
    always @ (*) begin
        if ((y <= 33) || (x >= 67 && y >= 34)) oled_data = 0;
        if (sw == 2'b00) begin // level 1
            // light blue
            if (pixel_index == 3501 || pixel_index == 3693 || pixel_index == 3885 || pixel_index == 3977 || pixel_index == 4169 || pixel_index == 4265 || pixel_index == 4360 || pixel_index == 4462 || pixel_index == 4557 || pixel_index == 4653 || pixel_index == 4750 || pixel_index == 5038 || pixel_index == 5133 || pixel_index == 5230 || pixel_index == 5416 || pixel_index == 5513 || pixel_index == 5608 || pixel_index == 5704 || pixel_index == 5801 || pixel_index == 3502 || pixel_index == 3597 || pixel_index == 3790 || pixel_index == 4072 || pixel_index == 4654 || pixel_index == 4845 || pixel_index == 4942 || pixel_index == 5325 || pixel_index == 5417 || pixel_index == 5800 || pixel_index == 3598 || pixel_index == 3694 || pixel_index == 3789 || pixel_index == 3886 || pixel_index == 3976 || pixel_index == 4073 || pixel_index == 4168 || pixel_index == 4558 || pixel_index == 4749 || pixel_index == 4846 || pixel_index == 4941 || pixel_index == 5037 || pixel_index == 5229 || pixel_index == 5326 || pixel_index == 5512 || pixel_index == 5705 || pixel_index == 4264 || pixel_index == 4361 || pixel_index == 4461 || pixel_index == 5134 || pixel_index == 5609) oled_data = 16'b0001111101111111;
            // white
            else if (((pixel_index >= 3503) && (pixel_index <= 3507)) || ((pixel_index >= 3599) && (pixel_index <= 3603)) || ((pixel_index >= 3695) && (pixel_index <= 3699)) || ((pixel_index >= 3791) && (pixel_index <= 3795)) || ((pixel_index >= 3887) && (pixel_index <= 3891)) || ((pixel_index >= 3978) && (pixel_index <= 3987)) || ((pixel_index >= 4074) && (pixel_index <= 4083)) || ((pixel_index >= 4170) && (pixel_index <= 4179)) || ((pixel_index >= 4266) && (pixel_index <= 4275)) || ((pixel_index >= 4362) && (pixel_index <= 4371)) || ((pixel_index >= 4463) && (pixel_index <= 4467)) || ((pixel_index >= 4559) && (pixel_index <= 4563)) || ((pixel_index >= 4655) && (pixel_index <= 4659)) || ((pixel_index >= 4751) && (pixel_index <= 4755)) || ((pixel_index >= 4847) && (pixel_index <= 4851)) || ((pixel_index >= 4943) && (pixel_index <= 4947)) || ((pixel_index >= 5039) && (pixel_index <= 5043)) || ((pixel_index >= 5135) && (pixel_index <= 5139)) || ((pixel_index >= 5231) && (pixel_index <= 5235)) || ((pixel_index >= 5327) && (pixel_index <= 5331)) || ((pixel_index >= 5418) && (pixel_index <= 5432)) || ((pixel_index >= 5514) && (pixel_index <= 5528)) || ((pixel_index >= 5610) && (pixel_index <= 5624)) || ((pixel_index >= 5706) && (pixel_index <= 5720)) || (pixel_index >= 5802) && (pixel_index <= 5816)) oled_data = 16'b1111111111111111;
            // pink
            else if (((pixel_index >= 3508) && (pixel_index <= 3509)) || ((pixel_index >= 3604) && (pixel_index <= 3605)) || pixel_index == 3700 || ((pixel_index >= 3796) && (pixel_index <= 3797)) || pixel_index == 3892 || ((pixel_index >= 3988) && (pixel_index <= 3989)) || pixel_index == 4084 || ((pixel_index >= 4180) && (pixel_index <= 4181)) || pixel_index == 4276 || ((pixel_index >= 4372) && (pixel_index <= 4373)) || pixel_index == 4468 || ((pixel_index >= 4564) && (pixel_index <= 4565)) || pixel_index == 4660 || ((pixel_index >= 4756) && (pixel_index <= 4757)) || pixel_index == 4852 || ((pixel_index >= 4948) && (pixel_index <= 4949)) || pixel_index == 5044 || ((pixel_index >= 5140) && (pixel_index <= 5141)) || pixel_index == 5237 || ((pixel_index >= 5332) && (pixel_index <= 5333)) || ((pixel_index >= 5433) && (pixel_index <= 5434)) || ((pixel_index >= 5529) && (pixel_index <= 5530)) || pixel_index == 5625 || ((pixel_index >= 5721) && (pixel_index <= 5722)) || pixel_index == 5818 || pixel_index == 3701 || pixel_index == 3893 || pixel_index == 4085 || pixel_index == 4277 || pixel_index == 4469 || pixel_index == 4661 || pixel_index == 4853 || pixel_index == 5045 || pixel_index == 5236 || pixel_index == 5626 || pixel_index == 5817) oled_data = 16'b1111100001011000;
            // bg
            else oled_data = 16'b0000000001000100;
        end
        if (sw[0] == 1) begin // level 2
            // light blue
            if (((pixel_index >= 3499) && (pixel_index <= 3500)) || ((pixel_index >= 3595) && (pixel_index <= 3596)) || pixel_index == 3691 || ((pixel_index >= 3787) && (pixel_index <= 3788)) || ((pixel_index >= 3883) && (pixel_index <= 3884)) || ((pixel_index >= 3974) && (pixel_index <= 3975)) || ((pixel_index >= 3989) && (pixel_index <= 3990)) || pixel_index == 4070 || pixel_index == 4086 || ((pixel_index >= 4166) && (pixel_index <= 4167)) || ((pixel_index >= 4181) && (pixel_index <= 4182)) || ((pixel_index >= 4262) && (pixel_index <= 4263)) || ((pixel_index >= 4277) && (pixel_index <= 4278)) || ((pixel_index >= 4358) && (pixel_index <= 4359)) || ((pixel_index >= 4373) && (pixel_index <= 4374)) || ((pixel_index >= 4464) && (pixel_index <= 4465)) || ((pixel_index >= 4560) && (pixel_index <= 4561)) || ((pixel_index >= 4656) && (pixel_index <= 4657)) || pixel_index == 4752 || ((pixel_index >= 4848) && (pixel_index <= 4849)) || ((pixel_index >= 4939) && (pixel_index <= 4940)) || ((pixel_index >= 5035) && (pixel_index <= 5036)) || pixel_index == 5131 || ((pixel_index >= 5227) && (pixel_index <= 5228)) || pixel_index == 5324 || ((pixel_index >= 5414) && (pixel_index <= 5415)) || pixel_index == 5511 || ((pixel_index >= 5606) && (pixel_index <= 5607)) || ((pixel_index >= 5702) && (pixel_index <= 5703)) || pixel_index == 5799 || pixel_index == 3692 || pixel_index == 4071 || pixel_index == 4085 || pixel_index == 4753 || pixel_index == 5132 || pixel_index == 5323 || pixel_index == 5510 || pixel_index == 5798) oled_data = 16'b0001011101111111;
            // white
            else if (((pixel_index >= 3501) && (pixel_index <= 3510)) || ((pixel_index >= 3597) && (pixel_index <= 3606)) || ((pixel_index >= 3693) && (pixel_index <= 3702)) || ((pixel_index >= 3789) && (pixel_index <= 3798)) || ((pixel_index >= 3885) && (pixel_index <= 3894)) || ((pixel_index >= 3976) && (pixel_index <= 3980)) || ((pixel_index >= 3991) && (pixel_index <= 3995)) || ((pixel_index >= 4072) && (pixel_index <= 4076)) || ((pixel_index >= 4087) && (pixel_index <= 4091)) || ((pixel_index >= 4168) && (pixel_index <= 4172)) || ((pixel_index >= 4183) && (pixel_index <= 4187)) || ((pixel_index >= 4264) && (pixel_index <= 4268)) || ((pixel_index >= 4279) && (pixel_index <= 4283)) || ((pixel_index >= 4360) && (pixel_index <= 4364)) || ((pixel_index >= 4375) && (pixel_index <= 4379)) || ((pixel_index >= 4466) && (pixel_index <= 4470)) || ((pixel_index >= 4562) && (pixel_index <= 4566)) || ((pixel_index >= 4658) && (pixel_index <= 4662)) || ((pixel_index >= 4754) && (pixel_index <= 4758)) || ((pixel_index >= 4850) && (pixel_index <= 4854)) || ((pixel_index >= 4941) && (pixel_index <= 4945)) || ((pixel_index >= 5037) && (pixel_index <= 5041)) || ((pixel_index >= 5133) && (pixel_index <= 5137)) || ((pixel_index >= 5229) && (pixel_index <= 5233)) || ((pixel_index >= 5325) && (pixel_index <= 5329)) || ((pixel_index >= 5416) && (pixel_index <= 5435)) || ((pixel_index >= 5512) && (pixel_index <= 5531)) || ((pixel_index >= 5608) && (pixel_index <= 5627)) || ((pixel_index >= 5704) && (pixel_index <= 5723)) || (pixel_index >= 5800) && (pixel_index <= 5819)) oled_data = 16'b1111111111111111;
            // pink
            else if (((pixel_index >= 3511) && (pixel_index <= 3512)) || ((pixel_index >= 3607) && (pixel_index <= 3608)) || pixel_index == 3703 || ((pixel_index >= 3799) && (pixel_index <= 3800)) || pixel_index == 3895 || ((pixel_index >= 3996) && (pixel_index <= 3997)) || ((pixel_index >= 4092) && (pixel_index <= 4093)) || pixel_index == 4188 || ((pixel_index >= 4284) && (pixel_index <= 4285)) || pixel_index == 4380 || pixel_index == 4471 || ((pixel_index >= 4567) && (pixel_index <= 4568)) || pixel_index == 4663 || ((pixel_index >= 4759) && (pixel_index <= 4760)) || pixel_index == 4855 || ((pixel_index >= 4946) && (pixel_index <= 4947)) || ((pixel_index >= 5042) && (pixel_index <= 5043)) || pixel_index == 5138 || pixel_index == 5234 || pixel_index == 5330 || pixel_index == 5436 || ((pixel_index >= 5532) && (pixel_index <= 5533)) || pixel_index == 5628 || ((pixel_index >= 5724) && (pixel_index <= 5725)) || pixel_index == 5821 || pixel_index == 3704 || pixel_index == 3896 || pixel_index == 4381 || pixel_index == 4664 || pixel_index == 4856 || pixel_index == 5139 || pixel_index == 5331 || pixel_index == 5437 || pixel_index == 5629 || pixel_index == 5820 || pixel_index == 4189 || pixel_index == 4472 || pixel_index == 5235) oled_data = 16'b1111100001011010;
            // bg
            else oled_data = 16'b0000000001000100;
        end
        if (sw[1] == 1) begin // level 3
            // light blue
            if (((pixel_index >= 3499) && (pixel_index <= 3500)) || ((pixel_index >= 3595) && (pixel_index <= 3596)) || pixel_index == 3691 || ((pixel_index >= 3787) && (pixel_index <= 3788)) || ((pixel_index >= 3883) && (pixel_index <= 3884)) || ((pixel_index >= 3974) && (pixel_index <= 3975)) || ((pixel_index >= 3989) && (pixel_index <= 3990)) || pixel_index == 4070 || pixel_index == 4086 || ((pixel_index >= 4166) && (pixel_index <= 4167)) || ((pixel_index >= 4181) && (pixel_index <= 4182)) || ((pixel_index >= 4262) && (pixel_index <= 4263)) || ((pixel_index >= 4277) && (pixel_index <= 4278)) || ((pixel_index >= 4358) && (pixel_index <= 4359)) || pixel_index == 4374 || ((pixel_index >= 4464) && (pixel_index <= 4465)) || ((pixel_index >= 4560) && (pixel_index <= 4561)) || ((pixel_index >= 4656) && (pixel_index <= 4657)) || pixel_index == 4752 || ((pixel_index >= 4848) && (pixel_index <= 4849)) || ((pixel_index >= 4934) && (pixel_index <= 4935)) || ((pixel_index >= 4949) && (pixel_index <= 4950)) || pixel_index == 5030 || ((pixel_index >= 5045) && (pixel_index <= 5046)) || ((pixel_index >= 5126) && (pixel_index <= 5127)) || pixel_index == 5141 || ((pixel_index >= 5222) && (pixel_index <= 5223)) || ((pixel_index >= 5237) && (pixel_index <= 5238)) || pixel_index == 5319 || ((pixel_index >= 5333) && (pixel_index <= 5334)) || ((pixel_index >= 5419) && (pixel_index <= 5420)) || pixel_index == 5515 || ((pixel_index >= 5611) && (pixel_index <= 5612)) || ((pixel_index >= 5707) && (pixel_index <= 5708)) || (pixel_index >= 5803) && (pixel_index <= 5804) || pixel_index == 3692 || pixel_index == 4071 || pixel_index == 4085 || pixel_index == 4373 || pixel_index == 4753 || pixel_index == 5031 || pixel_index == 5142 || pixel_index == 5318 || pixel_index == 5516) oled_data = 16'b0001011101111111;
            // white
            else if (((pixel_index >= 3501) && (pixel_index <= 3510)) || ((pixel_index >= 3597) && (pixel_index <= 3606)) || ((pixel_index >= 3693) && (pixel_index <= 3702)) || ((pixel_index >= 3789) && (pixel_index <= 3798)) || ((pixel_index >= 3885) && (pixel_index <= 3894)) || ((pixel_index >= 3976) && (pixel_index <= 3980)) || ((pixel_index >= 3991) && (pixel_index <= 3995)) || ((pixel_index >= 4072) && (pixel_index <= 4076)) || ((pixel_index >= 4087) && (pixel_index <= 4091)) || ((pixel_index >= 4168) && (pixel_index <= 4172)) || ((pixel_index >= 4183) && (pixel_index <= 4187)) || ((pixel_index >= 4264) && (pixel_index <= 4268)) || ((pixel_index >= 4279) && (pixel_index <= 4283)) || ((pixel_index >= 4360) && (pixel_index <= 4364)) || ((pixel_index >= 4375) && (pixel_index <= 4379)) || ((pixel_index >= 4466) && (pixel_index <= 4470)) || ((pixel_index >= 4562) && (pixel_index <= 4566)) || ((pixel_index >= 4658) && (pixel_index <= 4662)) || ((pixel_index >= 4754) && (pixel_index <= 4758)) || ((pixel_index >= 4850) && (pixel_index <= 4854)) || ((pixel_index >= 4936) && (pixel_index <= 4940)) || ((pixel_index >= 4951) && (pixel_index <= 4955)) || ((pixel_index >= 5032) && (pixel_index <= 5036)) || ((pixel_index >= 5047) && (pixel_index <= 5051)) || ((pixel_index >= 5128) && (pixel_index <= 5132)) || ((pixel_index >= 5143) && (pixel_index <= 5147)) || ((pixel_index >= 5224) && (pixel_index <= 5228)) || ((pixel_index >= 5239) && (pixel_index <= 5243)) || ((pixel_index >= 5320) && (pixel_index <= 5324)) || ((pixel_index >= 5335) && (pixel_index <= 5339)) || ((pixel_index >= 5421) && (pixel_index <= 5430)) || ((pixel_index >= 5517) && (pixel_index <= 5526)) || ((pixel_index >= 5613) && (pixel_index <= 5622)) || ((pixel_index >= 5709) && (pixel_index <= 5718)) || (pixel_index >= 5805) && (pixel_index <= 5814)) oled_data = 16'b1111111111111111;
            // pink
            else if (((pixel_index >= 3511) && (pixel_index <= 3512)) || pixel_index == 3607 || pixel_index == 3703 || ((pixel_index >= 3799) && (pixel_index <= 3800)) || pixel_index == 3896 || pixel_index == 3996 || ((pixel_index >= 4092) && (pixel_index <= 4093)) || pixel_index == 4189 || pixel_index == 4284 || pixel_index == 4380 || ((pixel_index >= 4471) && (pixel_index <= 4472)) || pixel_index == 4567 || ((pixel_index >= 4663) && (pixel_index <= 4664)) || pixel_index == 4760 || ((pixel_index >= 4855) && (pixel_index <= 4856)) || pixel_index == 4956 || pixel_index == 5053 || pixel_index == 5149 || ((pixel_index >= 5244) && (pixel_index <= 5245)) || pixel_index == 5340 || ((pixel_index >= 5431) && (pixel_index <= 5432)) || pixel_index == 5527 || pixel_index == 5623 || pixel_index == 5719 || pixel_index == 5816 || pixel_index == 3608 || pixel_index == 4568 || pixel_index == 5341 || pixel_index == 5528 || pixel_index == 3704 || pixel_index == 3895 || pixel_index == 3997 || pixel_index == 4188 || pixel_index == 4381 || pixel_index == 4759 || pixel_index == 4957 || pixel_index == 5148 || pixel_index == 5624 || pixel_index == 5720 || pixel_index == 5815 || pixel_index == 4285 || pixel_index == 5052) oled_data = 16'b1111100001011010;
            // bg
            else oled_data = 16'b0000000001000100;
        end
    end

endmodule

module comwait_data(input frame_rate, input sw, input [12:0] pixel_index, output reg [15:0] oled_data);
    reg [15:0] frame_count = 0;
    parameter picture_total_count = 8;
    
    wire [6:0] x = pixel_index % 96;
    wire [6:0] y = pixel_index / 96;
    
    always @ (posedge frame_rate) begin
        if (~sw) frame_count <= 0;
        else frame_count <= (frame_count == picture_total_count - 1) ? 0 : frame_count + 1;
    end
    
    always @ (*) begin
        if (y <= 33 || x <= 66) oled_data = 0;
        if (~sw) begin
            oled_data = 16'b0000000001000100;
        end
        else begin
            if (frame_count == 0) begin
                // white
                if (((pixel_index >= 3728) && (pixel_index <= 3729)) || ((pixel_index >= 3824) && (pixel_index <= 3825)) || ((pixel_index >= 3920) && (pixel_index <= 3921)) || ((pixel_index >= 4016) && (pixel_index <= 4017)) || ((pixel_index >= 4112) && (pixel_index <= 4113)) || ((pixel_index >= 4208) && (pixel_index <= 4209)) || ((pixel_index >= 4304) && (pixel_index <= 4305)) || (pixel_index >= 4400) && (pixel_index <= 4401)) oled_data = 16'b1111111111111111;
                // grey
                else if (pixel_index == 3912 || pixel_index == 3928 || pixel_index == 4008 || pixel_index == 4023 || pixel_index == 4025 || pixel_index == 4105 || pixel_index == 4107 || pixel_index == 4213 || pixel_index == 4215 || pixel_index == 4301 || pixel_index == 4308 || pixel_index == 4310 || pixel_index == 4397 || pixel_index == 4403 || pixel_index == 4405 || pixel_index == 4494 || pixel_index == 4678 || pixel_index == 4680 || pixel_index == 4699 || pixel_index == 4777 || pixel_index == 4779 || pixel_index == 4781 || pixel_index == 4788 || pixel_index == 4790 || pixel_index == 4794 || pixel_index == 4979 || pixel_index == 5070 || pixel_index == 5072 || pixel_index == 5163 || pixel_index == 5172 || pixel_index == 5174 || pixel_index == 5258 || pixel_index == 5260 || pixel_index == 5269 || pixel_index == 5271 || pixel_index == 5360 || pixel_index == 5367 || pixel_index == 5449 || pixel_index == 5464 || pixel_index == 5544 || pixel_index == 5552 || pixel_index == 3913 || pixel_index == 3929 || pixel_index == 4024 || pixel_index == 4106 || pixel_index == 4214 || pixel_index == 4309 || pixel_index == 4396 || pixel_index == 4404 || pixel_index == 4493 || pixel_index == 4679 || pixel_index == 4776 || pixel_index == 4778 || pixel_index == 4780 || pixel_index == 4789 || pixel_index == 4795 || pixel_index == 4980 || pixel_index == 5173 || pixel_index == 5259 || pixel_index == 5270 || pixel_index == 5361 || pixel_index == 5366 || pixel_index == 5368 || pixel_index == 5450 || pixel_index == 5463 || pixel_index == 5545 || pixel_index == 4009 || pixel_index == 4118 || pixel_index == 4120 || pixel_index == 4202 || pixel_index == 4204 || pixel_index == 4299 || pixel_index == 4398 || pixel_index == 4500 || pixel_index == 4682 || pixel_index == 4684 || pixel_index == 4693 || pixel_index == 4695 || pixel_index == 4697 || pixel_index == 4775 || pixel_index == 4791 || pixel_index == 4793 || pixel_index == 4974 || pixel_index == 5069 || pixel_index == 5073 || pixel_index == 5075 || pixel_index == 5077 || pixel_index == 5164 || pixel_index == 5168 || pixel_index == 5264 || pixel_index == 5353 || pixel_index == 5355 || pixel_index == 5448 || pixel_index == 5456 || pixel_index == 5553 || pixel_index == 5560 || pixel_index == 5648 || pixel_index == 5745 || pixel_index == 4010 || pixel_index == 4119 || pixel_index == 4203 || pixel_index == 4300 || pixel_index == 4499 || pixel_index == 4681 || pixel_index == 4683 || pixel_index == 4685 || pixel_index == 4692 || pixel_index == 4694 || pixel_index == 4696 || pixel_index == 4698 || pixel_index == 4774 || pixel_index == 4792 || pixel_index == 4973 || pixel_index == 5068 || pixel_index == 5076 || pixel_index == 5165 || pixel_index == 5169 || pixel_index == 5265 || pixel_index == 5354 || pixel_index == 5457 || pixel_index == 5465 || pixel_index == 5561 || pixel_index == 5649 || pixel_index == 5744) oled_data = 16'b1000010000010000;
                else oled_data = 16'b0000000001000100;
            end
            else if (frame_count == 1) begin
                // grey
                if (pixel_index == 3728 || pixel_index == 4010 || pixel_index == 4203 || pixel_index == 4300 || pixel_index == 4396 || pixel_index == 4693 || pixel_index == 4695 || pixel_index == 4697 || pixel_index == 4699 || pixel_index == 4774 || pixel_index == 4776 || pixel_index == 4778 || pixel_index == 4780 || pixel_index == 4792 || pixel_index == 4794 || pixel_index == 4973 || pixel_index == 5068 || pixel_index == 5070 || pixel_index == 5072 || pixel_index == 5077 || pixel_index == 5165 || pixel_index == 5173 || pixel_index == 5259 || pixel_index == 5264 || pixel_index == 5366 || pixel_index == 5368 || pixel_index == 5450 || pixel_index == 5545 || pixel_index == 5552 || pixel_index == 5561 || pixel_index == 5648 || pixel_index == 5745 || pixel_index == 3729 || pixel_index == 3825 || pixel_index == 3912 || pixel_index == 3920 || pixel_index == 4008 || pixel_index == 4016 || pixel_index == 4105 || pixel_index == 4107 || pixel_index == 4112 || pixel_index == 4208 || pixel_index == 4301 || pixel_index == 4305 || pixel_index == 4398 || pixel_index == 4400 || pixel_index == 4678 || pixel_index == 4680 || pixel_index == 4682 || pixel_index == 4684 || pixel_index == 4692 || pixel_index == 4790 || pixel_index == 4979 || pixel_index == 5073 || pixel_index == 5076 || pixel_index == 5163 || pixel_index == 5269 || pixel_index == 5271 || pixel_index == 5353 || pixel_index == 5361 || pixel_index == 5448 || pixel_index == 5456 || pixel_index == 5464 || pixel_index == 4009 || pixel_index == 4202 || pixel_index == 4204 || pixel_index == 4299 || pixel_index == 4397 || pixel_index == 4494 || pixel_index == 4694 || pixel_index == 4696 || pixel_index == 4698 || pixel_index == 4775 || pixel_index == 4777 || pixel_index == 4779 || pixel_index == 4781 || pixel_index == 4788 || pixel_index == 4791 || pixel_index == 4793 || pixel_index == 4795 || pixel_index == 4974 || pixel_index == 5069 || pixel_index == 5075 || pixel_index == 5164 || pixel_index == 5168 || pixel_index == 5172 || pixel_index == 5174 || pixel_index == 5258 || pixel_index == 5260 || pixel_index == 5265 || pixel_index == 5355 || pixel_index == 5367 || pixel_index == 5449 || pixel_index == 5544 || pixel_index == 5553 || pixel_index == 5560 || pixel_index == 5649 || pixel_index == 5744 || pixel_index == 3824 || pixel_index == 3913 || pixel_index == 3921 || pixel_index == 4017 || pixel_index == 4106 || pixel_index == 4113 || pixel_index == 4209 || pixel_index == 4304 || pixel_index == 4401 || pixel_index == 4493 || pixel_index == 4679 || pixel_index == 4681 || pixel_index == 4683 || pixel_index == 4685 || pixel_index == 4789 || pixel_index == 4980 || pixel_index == 5169 || pixel_index == 5270 || pixel_index == 5354 || pixel_index == 5360 || pixel_index == 5457 || pixel_index == 5463 || pixel_index == 5465) oled_data = 16'b1000010000010000;
                // white
                else if (((pixel_index >= 3928) && (pixel_index <= 3929)) || ((pixel_index >= 4023) && (pixel_index <= 4025)) || ((pixel_index >= 4118) && (pixel_index <= 4120)) || ((pixel_index >= 4213) && (pixel_index <= 4215)) || ((pixel_index >= 4308) && (pixel_index <= 4310)) || ((pixel_index >= 4403) && (pixel_index <= 4405)) || (pixel_index >= 4499) && (pixel_index <= 4500)) oled_data = 16'b1111111111111111;
                else oled_data = 16'b0000000001000100;
            end
            else if (frame_count == 2) begin
                // grey
                if (pixel_index == 3728 || pixel_index == 4010 || pixel_index == 4119 || pixel_index == 4203 || pixel_index == 4213 || pixel_index == 4300 || pixel_index == 4396 || pixel_index == 4403 || pixel_index == 4500 || pixel_index == 4774 || pixel_index == 4776 || pixel_index == 4778 || pixel_index == 4780 || pixel_index == 4973 || pixel_index == 5068 || pixel_index == 5070 || pixel_index == 5072 || pixel_index == 5165 || pixel_index == 5259 || pixel_index == 5264 || pixel_index == 5450 || pixel_index == 5465 || pixel_index == 5545 || pixel_index == 5552 || pixel_index == 5560 || pixel_index == 5648 || pixel_index == 5745 || pixel_index == 3729 || pixel_index == 3825 || pixel_index == 3912 || pixel_index == 3920 || pixel_index == 3928 || pixel_index == 4008 || pixel_index == 4016 || pixel_index == 4023 || pixel_index == 4025 || pixel_index == 4105 || pixel_index == 4107 || pixel_index == 4112 || pixel_index == 4208 || pixel_index == 4215 || pixel_index == 4301 || pixel_index == 4305 || pixel_index == 4309 || pixel_index == 4398 || pixel_index == 4400 || pixel_index == 4678 || pixel_index == 4680 || pixel_index == 4682 || pixel_index == 4684 || pixel_index == 4979 || pixel_index == 5073 || pixel_index == 5076 || pixel_index == 5163 || pixel_index == 5172 || pixel_index == 5174 || pixel_index == 5269 || pixel_index == 5271 || pixel_index == 5353 || pixel_index == 5361 || pixel_index == 5367 || pixel_index == 5448 || pixel_index == 5456 || pixel_index == 5464 || pixel_index == 3824 || pixel_index == 3913 || pixel_index == 3921 || pixel_index == 3929 || pixel_index == 4017 || pixel_index == 4024 || pixel_index == 4106 || pixel_index == 4113 || pixel_index == 4209 || pixel_index == 4304 || pixel_index == 4310 || pixel_index == 4401 || pixel_index == 4405 || pixel_index == 4493 || pixel_index == 4679 || pixel_index == 4681 || pixel_index == 4683 || pixel_index == 4685 || pixel_index == 4980 || pixel_index == 5077 || pixel_index == 5169 || pixel_index == 5173 || pixel_index == 5270 || pixel_index == 5354 || pixel_index == 5360 || pixel_index == 5366 || pixel_index == 5457 || pixel_index == 5463 || pixel_index == 4009 || pixel_index == 4118 || pixel_index == 4120 || pixel_index == 4202 || pixel_index == 4204 || pixel_index == 4214 || pixel_index == 4299 || pixel_index == 4308 || pixel_index == 4397 || pixel_index == 4404 || pixel_index == 4494 || pixel_index == 4499 || pixel_index == 4775 || pixel_index == 4777 || pixel_index == 4779 || pixel_index == 4781 || pixel_index == 4974 || pixel_index == 5069 || pixel_index == 5075 || pixel_index == 5164 || pixel_index == 5168 || pixel_index == 5258 || pixel_index == 5260 || pixel_index == 5265 || pixel_index == 5355 || pixel_index == 5368 || pixel_index == 5449 || pixel_index == 5544 || pixel_index == 5553 || pixel_index == 5561 || pixel_index == 5649 || pixel_index == 5744) oled_data = 16'b1000010000010000;
                // white
                else if (((pixel_index >= 4692) && (pixel_index <= 4699)) || (pixel_index >= 4788) && (pixel_index <= 4795)) oled_data = 16'b1111111111111111;
                else oled_data = 16'b0000000001000100;
            end
            else if (frame_count == 3) begin
                // grey
                if (pixel_index == 3728 || pixel_index == 4010 || pixel_index == 4119 || pixel_index == 4203 || pixel_index == 4213 || pixel_index == 4300 || pixel_index == 4396 || pixel_index == 4403 || pixel_index == 4500 || pixel_index == 4693 || pixel_index == 4695 || pixel_index == 4774 || pixel_index == 4776 || pixel_index == 4778 || pixel_index == 4780 || pixel_index == 4790 || pixel_index == 4792 || pixel_index == 4794 || pixel_index == 4973 || pixel_index == 5068 || pixel_index == 5070 || pixel_index == 5072 || pixel_index == 5165 || pixel_index == 5259 || pixel_index == 5264 || pixel_index == 5450 || pixel_index == 5545 || pixel_index == 5552 || pixel_index == 5648 || pixel_index == 5745 || pixel_index == 3729 || pixel_index == 3825 || pixel_index == 3912 || pixel_index == 3920 || pixel_index == 3928 || pixel_index == 4008 || pixel_index == 4016 || pixel_index == 4023 || pixel_index == 4025 || pixel_index == 4105 || pixel_index == 4107 || pixel_index == 4112 || pixel_index == 4208 || pixel_index == 4215 || pixel_index == 4301 || pixel_index == 4305 || pixel_index == 4309 || pixel_index == 4398 || pixel_index == 4400 || pixel_index == 4678 || pixel_index == 4680 || pixel_index == 4682 || pixel_index == 4684 || pixel_index == 4692 || pixel_index == 4696 || pixel_index == 4698 || pixel_index == 5073 || pixel_index == 5163 || pixel_index == 5353 || pixel_index == 5361 || pixel_index == 5448 || pixel_index == 5456 || pixel_index == 3824 || pixel_index == 3913 || pixel_index == 3921 || pixel_index == 3929 || pixel_index == 4017 || pixel_index == 4024 || pixel_index == 4106 || pixel_index == 4113 || pixel_index == 4209 || pixel_index == 4304 || pixel_index == 4310 || pixel_index == 4401 || pixel_index == 4405 || pixel_index == 4493 || pixel_index == 4679 || pixel_index == 4681 || pixel_index == 4683 || pixel_index == 4685 || pixel_index == 4697 || pixel_index == 4699 || pixel_index == 4788 || pixel_index == 5169 || pixel_index == 5354 || pixel_index == 5360 || pixel_index == 5457 || pixel_index == 4009 || pixel_index == 4118 || pixel_index == 4120 || pixel_index == 4202 || pixel_index == 4204 || pixel_index == 4214 || pixel_index == 4299 || pixel_index == 4308 || pixel_index == 4397 || pixel_index == 4404 || pixel_index == 4494 || pixel_index == 4499 || pixel_index == 4694 || pixel_index == 4775 || pixel_index == 4777 || pixel_index == 4779 || pixel_index == 4781 || pixel_index == 4789 || pixel_index == 4791 || pixel_index == 4793 || pixel_index == 4795 || pixel_index == 4974 || pixel_index == 5069 || pixel_index == 5164 || pixel_index == 5168 || pixel_index == 5258 || pixel_index == 5260 || pixel_index == 5265 || pixel_index == 5355 || pixel_index == 5449 || pixel_index == 5544 || pixel_index == 5553 || pixel_index == 5649 || pixel_index == 5744) oled_data = 16'b1000010000010000;
                // white
                else if (((pixel_index >= 4979) && (pixel_index <= 4980)) || ((pixel_index >= 5075) && (pixel_index <= 5077)) || ((pixel_index >= 5172) && (pixel_index <= 5174)) || ((pixel_index >= 5269) && (pixel_index <= 5271)) || ((pixel_index >= 5366) && (pixel_index <= 5368)) || ((pixel_index >= 5463) && (pixel_index <= 5465)) || (pixel_index >= 5560) && (pixel_index <= 5561)) oled_data = 16'b1111111111111111;
                else oled_data = 16'b0000000001000100;
            end
            else if (frame_count == 4) begin
                // grey
                if (pixel_index == 3728 || pixel_index == 4010 || pixel_index == 4119 || pixel_index == 4203 || pixel_index == 4213 || pixel_index == 4300 || pixel_index == 4396 || pixel_index == 4403 || pixel_index == 4500 || pixel_index == 4693 || pixel_index == 4695 || pixel_index == 4774 || pixel_index == 4776 || pixel_index == 4778 || pixel_index == 4780 || pixel_index == 4790 || pixel_index == 4792 || pixel_index == 4794 || pixel_index == 4973 || pixel_index == 5068 || pixel_index == 5070 || pixel_index == 5075 || pixel_index == 5077 || pixel_index == 5165 || pixel_index == 5172 || pixel_index == 5259 || pixel_index == 5450 || pixel_index == 5545 || pixel_index == 3729 || pixel_index == 3825 || pixel_index == 3912 || pixel_index == 3920 || pixel_index == 3928 || pixel_index == 4008 || pixel_index == 4016 || pixel_index == 4023 || pixel_index == 4025 || pixel_index == 4105 || pixel_index == 4107 || pixel_index == 4112 || pixel_index == 4208 || pixel_index == 4215 || pixel_index == 4301 || pixel_index == 4305 || pixel_index == 4309 || pixel_index == 4398 || pixel_index == 4400 || pixel_index == 4678 || pixel_index == 4680 || pixel_index == 4682 || pixel_index == 4684 || pixel_index == 4692 || pixel_index == 4696 || pixel_index == 4698 || pixel_index == 4979 || pixel_index == 5163 || pixel_index == 5174 || pixel_index == 5270 || pixel_index == 5353 || pixel_index == 5366 || pixel_index == 5368 || pixel_index == 5448 || pixel_index == 5463 || pixel_index == 5465 || pixel_index == 5561 || pixel_index == 3824 || pixel_index == 3913 || pixel_index == 3921 || pixel_index == 3929 || pixel_index == 4017 || pixel_index == 4024 || pixel_index == 4106 || pixel_index == 4113 || pixel_index == 4209 || pixel_index == 4304 || pixel_index == 4310 || pixel_index == 4401 || pixel_index == 4405 || pixel_index == 4493 || pixel_index == 4679 || pixel_index == 4681 || pixel_index == 4683 || pixel_index == 4685 || pixel_index == 4697 || pixel_index == 4699 || pixel_index == 4788 || pixel_index == 4980 || pixel_index == 5269 || pixel_index == 5271 || pixel_index == 5354 || pixel_index == 5367 || pixel_index == 5464 || pixel_index == 5560 || pixel_index == 4009 || pixel_index == 4118 || pixel_index == 4120 || pixel_index == 4202 || pixel_index == 4204 || pixel_index == 4214 || pixel_index == 4299 || pixel_index == 4308 || pixel_index == 4397 || pixel_index == 4404 || pixel_index == 4494 || pixel_index == 4499 || pixel_index == 4694 || pixel_index == 4775 || pixel_index == 4777 || pixel_index == 4779 || pixel_index == 4781 || pixel_index == 4789 || pixel_index == 4791 || pixel_index == 4793 || pixel_index == 4795 || pixel_index == 4974 || pixel_index == 5069 || pixel_index == 5076 || pixel_index == 5164 || pixel_index == 5173 || pixel_index == 5258 || pixel_index == 5260 || pixel_index == 5355 || pixel_index == 5449 || pixel_index == 5544) oled_data = 16'b1000010000010000;
                // white
                else if (((pixel_index >= 5072) && (pixel_index <= 5073)) || ((pixel_index >= 5168) && (pixel_index <= 5169)) || ((pixel_index >= 5264) && (pixel_index <= 5265)) || ((pixel_index >= 5360) && (pixel_index <= 5361)) || ((pixel_index >= 5456) && (pixel_index <= 5457)) || ((pixel_index >= 5552) && (pixel_index <= 5553)) || ((pixel_index >= 5648) && (pixel_index <= 5649)) || (pixel_index >= 5744) && (pixel_index <= 5745)) oled_data = 16'b1111111111111111;
                else oled_data = 16'b0000000001000100;
            end
            else if (frame_count == 5) begin
                // grey
                if (pixel_index == 3728 || pixel_index == 4010 || pixel_index == 4119 || pixel_index == 4203 || pixel_index == 4213 || pixel_index == 4300 || pixel_index == 4396 || pixel_index == 4403 || pixel_index == 4500 || pixel_index == 4693 || pixel_index == 4695 || pixel_index == 4774 || pixel_index == 4776 || pixel_index == 4778 || pixel_index == 4780 || pixel_index == 4790 || pixel_index == 4792 || pixel_index == 4794 || pixel_index == 5073 || pixel_index == 5077 || pixel_index == 5173 || pixel_index == 5265 || pixel_index == 5271 || pixel_index == 5360 || pixel_index == 5457 || pixel_index == 5465 || pixel_index == 5648 || pixel_index == 3729 || pixel_index == 3825 || pixel_index == 3912 || pixel_index == 3920 || pixel_index == 3928 || pixel_index == 4008 || pixel_index == 4016 || pixel_index == 4023 || pixel_index == 4025 || pixel_index == 4105 || pixel_index == 4107 || pixel_index == 4112 || pixel_index == 4208 || pixel_index == 4215 || pixel_index == 4301 || pixel_index == 4305 || pixel_index == 4309 || pixel_index == 4398 || pixel_index == 4400 || pixel_index == 4678 || pixel_index == 4680 || pixel_index == 4682 || pixel_index == 4684 || pixel_index == 4692 || pixel_index == 4696 || pixel_index == 4698 || pixel_index == 4979 || pixel_index == 5072 || pixel_index == 5076 || pixel_index == 5264 || pixel_index == 5270 || pixel_index == 5367 || pixel_index == 5463 || pixel_index == 5552 || pixel_index == 5561 || pixel_index == 5745 || pixel_index == 3824 || pixel_index == 3913 || pixel_index == 3921 || pixel_index == 3929 || pixel_index == 4017 || pixel_index == 4024 || pixel_index == 4106 || pixel_index == 4113 || pixel_index == 4209 || pixel_index == 4304 || pixel_index == 4310 || pixel_index == 4401 || pixel_index == 4405 || pixel_index == 4493 || pixel_index == 4679 || pixel_index == 4681 || pixel_index == 4683 || pixel_index == 4685 || pixel_index == 4697 || pixel_index == 4699 || pixel_index == 4788 || pixel_index == 4980 || pixel_index == 5075 || pixel_index == 5269 || pixel_index == 5366 || pixel_index == 5368 || pixel_index == 5553 || pixel_index == 5560 || pixel_index == 4009 || pixel_index == 4118 || pixel_index == 4120 || pixel_index == 4202 || pixel_index == 4204 || pixel_index == 4214 || pixel_index == 4299 || pixel_index == 4308 || pixel_index == 4397 || pixel_index == 4404 || pixel_index == 4494 || pixel_index == 4499 || pixel_index == 4694 || pixel_index == 4775 || pixel_index == 4777 || pixel_index == 4779 || pixel_index == 4781 || pixel_index == 4789 || pixel_index == 4791 || pixel_index == 4793 || pixel_index == 4795 || ((pixel_index >= 5168) && (pixel_index <= 5169)) || pixel_index == 5172 || pixel_index == 5174 || pixel_index == 5361 || pixel_index == 5456 || pixel_index == 5464 || pixel_index == 5649 || pixel_index == 5744) oled_data = 16'b1000010000010000;
                // white
                else if (((pixel_index >= 4973) && (pixel_index <= 4974)) || ((pixel_index >= 5068) && (pixel_index <= 5070)) || ((pixel_index >= 5163) && (pixel_index <= 5165)) || ((pixel_index >= 5258) && (pixel_index <= 5260)) || ((pixel_index >= 5353) && (pixel_index <= 5355)) || ((pixel_index >= 5448) && (pixel_index <= 5450)) || (pixel_index >= 5544) && (pixel_index <= 5545)) oled_data = 16'b1111111111111111;
                else oled_data = 16'b0000000001000100;
            end
            else if (frame_count == 6) begin
                // grey
                if (pixel_index == 3728 || pixel_index == 4010 || pixel_index == 4119 || pixel_index == 4203 || pixel_index == 4213 || pixel_index == 4300 || pixel_index == 4396 || pixel_index == 4403 || pixel_index == 4500 || pixel_index == 4692 || pixel_index == 4696 || pixel_index == 4698 || pixel_index == 4789 || pixel_index == 4791 || pixel_index == 4793 || pixel_index == 4795 || pixel_index == 4973 || pixel_index == 4979 || pixel_index == 5072 || pixel_index == 5163 || pixel_index == 5165 || pixel_index == 5173 || pixel_index == 5258 || pixel_index == 5260 || pixel_index == 5360 || pixel_index == 5366 || pixel_index == 5368 || pixel_index == 5457 || pixel_index == 5465 || pixel_index == 5552 || pixel_index == 5561 || pixel_index == 3729 || pixel_index == 3825 || pixel_index == 3912 || pixel_index == 3920 || pixel_index == 3928 || pixel_index == 4008 || pixel_index == 4016 || pixel_index == 4023 || pixel_index == 4025 || pixel_index == 4105 || pixel_index == 4107 || pixel_index == 4112 || pixel_index == 4208 || pixel_index == 4215 || pixel_index == 4301 || pixel_index == 4305 || pixel_index == 4309 || pixel_index == 4398 || pixel_index == 4400 || pixel_index == 4693 || pixel_index == 4695 || pixel_index == 4974 || pixel_index == 4980 || pixel_index == 5068 || pixel_index == 5077 || pixel_index == 5168 || pixel_index == 5265 || pixel_index == 5270 || pixel_index == 5353 || pixel_index == 5355 || pixel_index == 5448 || pixel_index == 5450 || pixel_index == 5463 || pixel_index == 5545 || pixel_index == 5649 || pixel_index == 5744 || pixel_index == 3824 || pixel_index == 3913 || pixel_index == 3921 || pixel_index == 3929 || pixel_index == 4017 || pixel_index == 4024 || pixel_index == 4106 || pixel_index == 4113 || pixel_index == 4209 || pixel_index == 4304 || pixel_index == 4310 || pixel_index == 4401 || pixel_index == 4405 || pixel_index == 4493 || pixel_index == 4694 || pixel_index == 5069 || pixel_index == 5076 || pixel_index == 5264 || pixel_index == 5271 || pixel_index == 5354 || pixel_index == 5449 || pixel_index == 5648 || pixel_index == 5745 || pixel_index == 4009 || pixel_index == 4118 || pixel_index == 4120 || pixel_index == 4202 || pixel_index == 4204 || pixel_index == 4214 || pixel_index == 4299 || pixel_index == 4308 || pixel_index == 4397 || pixel_index == 4404 || pixel_index == 4494 || pixel_index == 4499 || pixel_index == 4697 || pixel_index == 4699 || pixel_index == 4788 || pixel_index == 4790 || pixel_index == 4792 || pixel_index == 4794 || pixel_index == 5070 || pixel_index == 5073 || pixel_index == 5075 || pixel_index == 5164 || pixel_index == 5169 || pixel_index == 5172 || pixel_index == 5174 || pixel_index == 5259 || pixel_index == 5269 || pixel_index == 5361 || pixel_index == 5367 || pixel_index == 5456 || pixel_index == 5464 || pixel_index == 5544 || pixel_index == 5553 || pixel_index == 5560) oled_data = 16'b1000010000010000;
                // white
                else if (((pixel_index >= 4678) && (pixel_index <= 4685)) || (pixel_index >= 4774) && (pixel_index <= 4781)) oled_data = 16'b1111111111111111;
                else oled_data = 16'b0000000001000100;
            end
            else if (frame_count == 7) begin
                // grey
                if (pixel_index == 3728 || pixel_index == 3920 || pixel_index == 3928 || pixel_index == 4023 || pixel_index == 4025 || pixel_index == 4113 || pixel_index == 4119 || pixel_index == 4208 || pixel_index == 4500 || pixel_index == 4681 || pixel_index == 4683 || pixel_index == 4685 || pixel_index == 4698 || pixel_index == 4973 || pixel_index == 4979 || pixel_index == 5068 || pixel_index == 5072 || pixel_index == 5163 || pixel_index == 5174 || pixel_index == 5360 || pixel_index == 5368 || pixel_index == 5448 || pixel_index == 5545 || pixel_index == 5648 || pixel_index == 5745 || pixel_index == 3729 || pixel_index == 3825 || pixel_index == 4016 || pixel_index == 4213 || pixel_index == 4215 || pixel_index == 4304 || pixel_index == 4308 || pixel_index == 4310 || pixel_index == 4401 || pixel_index == 4403 || pixel_index == 4405 || pixel_index == 4678 || pixel_index == 4680 || pixel_index == 4684 || pixel_index == 4692 || pixel_index == 4694 || pixel_index == 4696 || pixel_index == 4699 || pixel_index == 4774 || pixel_index == 4777 || pixel_index == 4779 || pixel_index == 4788 || pixel_index == 4791 || pixel_index == 4793 || pixel_index == 4974 || pixel_index == 5075 || pixel_index == 5077 || pixel_index == 5165 || pixel_index == 5168 || pixel_index == 5172 || pixel_index == 5259 || pixel_index == 5265 || pixel_index == 5270 || pixel_index == 5353 || pixel_index == 5367 || pixel_index == 5450 || pixel_index == 5456 || pixel_index == 5464 || pixel_index == 5552 || pixel_index == 5561 || pixel_index == 3824 || pixel_index == 4017 || pixel_index == 4214 || pixel_index == 4305 || pixel_index == 4309 || pixel_index == 4400 || pixel_index == 4404 || pixel_index == 4679 || pixel_index == 4693 || pixel_index == 4695 || pixel_index == 4775 || pixel_index == 4778 || pixel_index == 4780 || pixel_index == 4789 || pixel_index == 4792 || pixel_index == 4794 || pixel_index == 5070 || pixel_index == 5076 || pixel_index == 5169 || pixel_index == 5258 || pixel_index == 5260 || pixel_index == 5264 || pixel_index == 5269 || pixel_index == 5271 || pixel_index == 5354 || pixel_index == 5366 || pixel_index == 5457 || pixel_index == 5465 || pixel_index == 5553 || pixel_index == 5560 || pixel_index == 3921 || pixel_index == 3929 || pixel_index == 4024 || pixel_index == 4112 || pixel_index == 4118 || pixel_index == 4120 || pixel_index == 4209 || pixel_index == 4499 || pixel_index == 4682 || pixel_index == 4697 || pixel_index == 4776 || pixel_index == 4781 || pixel_index == 4790 || pixel_index == 4795 || pixel_index == 4980 || pixel_index == 5069 || pixel_index == 5073 || pixel_index == 5164 || pixel_index == 5173 || pixel_index == 5355 || pixel_index == 5361 || pixel_index == 5449 || pixel_index == 5463 || pixel_index == 5544 || pixel_index == 5649 || pixel_index == 5744) oled_data = 16'b1000010000010000;
                // white
                else if (((pixel_index >= 3912) && (pixel_index <= 3913)) || ((pixel_index >= 4008) && (pixel_index <= 4010)) || ((pixel_index >= 4105) && (pixel_index <= 4107)) || ((pixel_index >= 4202) && (pixel_index <= 4204)) || ((pixel_index >= 4299) && (pixel_index <= 4301)) || ((pixel_index >= 4396) && (pixel_index <= 4398)) || (pixel_index >= 4493) && (pixel_index <= 4494)) oled_data = 16'b1111111111111111;
                else oled_data = 16'b0000000001000100;
            end
        end
    end

endmodule