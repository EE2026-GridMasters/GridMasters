`timescale 1ns / 1ps

module display_home_page(
    input [12:0] pixel_index,
    output reg [15:0] oled_data
    );
    
    parameter PINK_HEX = 16'hF899;
    parameter BLUE_HEX = 16'h177F;
    parameter BG_BLUE_HEX = 16'b0000000001000100;
    parameter WHITE_HEX = 16'hFFFF;
    
    always @(*) begin
        if ((pixel_index >= 1365 && pixel_index <= 1367) || (pixel_index >= 1390 && pixel_index <= 1392) || (pixel_index >= 1407 && pixel_index <= 1409) || (pixel_index >= 1428 && pixel_index <= 1430) || (pixel_index >= 1461 && pixel_index <= 1463) || (pixel_index >= 1486 && pixel_index <= 1488) || (pixel_index >= 1503 && pixel_index <= 1505) || (pixel_index >= 1524 && pixel_index <= 1526) || (pixel_index >= 1557 && pixel_index <= 1559) || (pixel_index >= 1582 && pixel_index <= 1584) || (pixel_index >= 1599 && pixel_index <= 1601) || (pixel_index >= 1620 && pixel_index <= 1622) || (pixel_index >= 1653 && pixel_index <= 1655) || (pixel_index >= 1678 && pixel_index <= 1680) || (pixel_index >= 1695 && pixel_index <= 1697) || (pixel_index >= 1716 && pixel_index <= 1718) || (pixel_index >= 1749 && pixel_index <= 1751) || (pixel_index >= 1774 && pixel_index <= 1776) || (pixel_index >= 1791 && pixel_index <= 1793) || (pixel_index >= 1812 && pixel_index <= 1814) || (pixel_index >= 1836 && pixel_index <= 1838) || (pixel_index >= 1849 && pixel_index <= 1851) || (pixel_index >= 1861 && pixel_index <= 1863) || (pixel_index >= 1875 && pixel_index <= 1877) || (pixel_index >= 1887 && pixel_index <= 1889) || (pixel_index >= 1899 && pixel_index <= 1901) || (pixel_index >= 1913 && pixel_index <= 1915) || (pixel_index >= 1932 && pixel_index <= 1934) || (pixel_index >= 1945 && pixel_index <= 1947) || (pixel_index >= 1957 && pixel_index <= 1959) || (pixel_index >= 1971 && pixel_index <= 1973) || (pixel_index >= 1983 && pixel_index <= 1985) || (pixel_index >= 1995 && pixel_index <= 1997) || (pixel_index >= 2009 && pixel_index <= 2011) || (pixel_index >= 2028 && pixel_index <= 2030) || (pixel_index >= 2041 && pixel_index <= 2043) || (pixel_index >= 2053 && pixel_index <= 2055) || (pixel_index >= 2067 && pixel_index <= 2069) || (pixel_index >= 2079 && pixel_index <= 2081) || (pixel_index >= 2091 && pixel_index <= 2093) || (pixel_index >= 2105 && pixel_index <= 2107) || (pixel_index >= 2124 && pixel_index <= 2126) || (pixel_index >= 2137 && pixel_index <= 2139) || (pixel_index >= 2149 && pixel_index <= 2151) || (pixel_index >= 2163 && pixel_index <= 2165) || (pixel_index >= 2175 && pixel_index <= 2177) || (pixel_index >= 2187 && pixel_index <= 2189) || (pixel_index >= 2201 && pixel_index <= 2203) || (pixel_index >= 2220 && pixel_index <= 2222) || (pixel_index >= 2233 && pixel_index <= 2235) || (pixel_index >= 2245 && pixel_index <= 2247) || (pixel_index >= 2259 && pixel_index <= 2261) || (pixel_index >= 2271 && pixel_index <= 2273) || (pixel_index >= 2283 && pixel_index <= 2285) || (pixel_index >= 2297 && pixel_index <= 2299) || (pixel_index >= 2316 && pixel_index <= 2318) || (pixel_index >= 2341 && pixel_index <= 2343) || (pixel_index >= 2355 && pixel_index <= 2357) || (pixel_index >= 2367 && pixel_index <= 2369) || (pixel_index >= 2379 && pixel_index <= 2381) || (pixel_index >= 2393 && pixel_index <= 2395) || (pixel_index >= 2412 && pixel_index <= 2414) || (pixel_index >= 2451 && pixel_index <= 2453) || (pixel_index >= 2463 && pixel_index <= 2465) || (pixel_index >= 2475 && pixel_index <= 2477) || (pixel_index >= 2489 && pixel_index <= 2491) || (pixel_index >= 2508 && pixel_index <= 2510) || (pixel_index >= 2543 && pixel_index <= 2545) || (pixel_index >= 2559 && pixel_index <= 2561) || (pixel_index >= 2571 && pixel_index <= 2573) || (pixel_index >= 2585 && pixel_index <= 2587) || (pixel_index >= 2604 && pixel_index <= 2605) || (pixel_index >= 2617 && pixel_index <= 2619) || (pixel_index >= 2639 && pixel_index <= 2641) || (pixel_index >= 2655 && pixel_index <= 2657) || (pixel_index >= 2667 && pixel_index <= 2669) || (pixel_index >= 2681 && pixel_index <= 2683) || (pixel_index >= 2700 && pixel_index <= 2701) || (pixel_index >= 2713 && pixel_index <= 2715) || (pixel_index >= 2735 && pixel_index <= 2737) || (pixel_index >= 2751 && pixel_index <= 2753) || (pixel_index >= 2763 && pixel_index <= 2765) || (pixel_index >= 2777 && pixel_index <= 2779) || (pixel_index >= 2796 && pixel_index <= 2797) || (pixel_index >= 2809 && pixel_index <= 2811) || (pixel_index >= 2835 && pixel_index <= 2837) || (pixel_index >= 2847 && pixel_index <= 2849) || (pixel_index >= 2859 && pixel_index <= 2861) || (pixel_index >= 2873 && pixel_index <= 2875) || (pixel_index >= 2892 && pixel_index <= 2893) || (pixel_index >= 2905 && pixel_index <= 2907) || (pixel_index >= 2917 && pixel_index <= 2919) || (pixel_index >= 2931 && pixel_index <= 2933) || (pixel_index >= 2943 && pixel_index <= 2945) || (pixel_index >= 2955 && pixel_index <= 2957) || (pixel_index >= 2969 && pixel_index <= 2971) || (pixel_index >= 2988 && pixel_index <= 2989) || (pixel_index >= 3001 && pixel_index <= 3003) || (pixel_index >= 3013 && pixel_index <= 3015) || (pixel_index >= 3027 && pixel_index <= 3029) || (pixel_index >= 3039 && pixel_index <= 3041) || (pixel_index >= 3051 && pixel_index <= 3053) || (pixel_index >= 3065 && pixel_index <= 3067) || (pixel_index >= 3084 && pixel_index <= 3086) || (pixel_index >= 3097 && pixel_index <= 3099) || (pixel_index >= 3109 && pixel_index <= 3111) || (pixel_index >= 3123 && pixel_index <= 3125) || (pixel_index >= 3135 && pixel_index <= 3137) || (pixel_index >= 3147 && pixel_index <= 3149) || (pixel_index >= 3161 && pixel_index <= 3163) || (pixel_index >= 3180 && pixel_index <= 3182) || (pixel_index >= 3193 && pixel_index <= 3195) || (pixel_index >= 3205 && pixel_index <= 3207) || (pixel_index >= 3219 && pixel_index <= 3221) || (pixel_index >= 3231 && pixel_index <= 3233) || (pixel_index >= 3243 && pixel_index <= 3245) || (pixel_index >= 3257 && pixel_index <= 3259) || (pixel_index >= 3276 && pixel_index <= 3278) || (pixel_index >= 3289 && pixel_index <= 3291) || (pixel_index >= 3301 && pixel_index <= 3303) || (pixel_index >= 3315 && pixel_index <= 3317) || (pixel_index >= 3327 && pixel_index <= 3329) || (pixel_index >= 3339 && pixel_index <= 3341) || (pixel_index >= 3353 && pixel_index <= 3355) || (pixel_index >= 3372 && pixel_index <= 3374) || (pixel_index >= 3385 && pixel_index <= 3387) || (pixel_index >= 3397 && pixel_index <= 3399) || (pixel_index >= 3411 && pixel_index <= 3413) || (pixel_index >= 3423 && pixel_index <= 3425) || (pixel_index >= 3435 && pixel_index <= 3437) || (pixel_index >= 3449 && pixel_index <= 3451) || (pixel_index >= 3477 && pixel_index <= 3479) || (pixel_index >= 3493 && pixel_index <= 3495) || (pixel_index >= 3507 && pixel_index <= 3509) || (pixel_index >= 3519 && pixel_index <= 3521) || (pixel_index >= 3540 && pixel_index <= 3542) || (pixel_index >= 3573 && pixel_index <= 3575) || (pixel_index >= 3589 && pixel_index <= 3591) || (pixel_index >= 3603 && pixel_index <= 3605) || (pixel_index >= 3615 && pixel_index <= 3617) || (pixel_index >= 3636 && pixel_index <= 3638) || (pixel_index >= 3669 && pixel_index <= 3671) || (pixel_index >= 3685 && pixel_index <= 3687) || (pixel_index >= 3699 && pixel_index <= 3701) || (pixel_index >= 3711 && pixel_index <= 3713) || (pixel_index >= 3732 && pixel_index <= 3734) || (pixel_index >= 3765 && pixel_index <= 3767) || (pixel_index >= 3781 && pixel_index <= 3783) || (pixel_index >= 3795 && pixel_index <= 3797) || (pixel_index >= 3807 && pixel_index <= 3809) || (pixel_index >= 3828 && pixel_index <= 3830) || (pixel_index >= 3861 && pixel_index <= 3863) || (pixel_index >= 3877 && pixel_index <= 3879) || (pixel_index >= 3891 && pixel_index <= 3893) || (pixel_index >= 3903 && pixel_index <= 3905) || (pixel_index >= 3924 && pixel_index <= 3926)) begin
            oled_data = PINK_HEX;
        end else if ((pixel_index >= 1353 && pixel_index <= 1355) || (pixel_index >= 1374 && pixel_index <= 1376) || (pixel_index >= 1400 && pixel_index <= 1402) || (pixel_index >= 1412 && pixel_index <= 1414) || (pixel_index >= 1449 && pixel_index <= 1450) || (pixel_index >= 1470 && pixel_index <= 1472) || (pixel_index >= 1496 && pixel_index <= 1497) || (pixel_index >= 1508 && pixel_index <= 1509) || (pixel_index >= 1545 && pixel_index <= 1546) || (pixel_index >= 1566 && pixel_index <= 1568) || (pixel_index >= 1592 && pixel_index <= 1593) || (pixel_index >= 1604 && pixel_index <= 1605) || (pixel_index >= 1641 && pixel_index <= 1642) || (pixel_index >= 1662 && pixel_index <= 1664) || (pixel_index >= 1688 && pixel_index <= 1689) || (pixel_index >= 1700 && pixel_index <= 1701) || (pixel_index >= 1737 && pixel_index <= 1739) || (pixel_index >= 1758 && pixel_index <= 1760) || (pixel_index >= 1784 && pixel_index <= 1785) || (pixel_index >= 1796 && pixel_index <= 1797) || (pixel_index >= 1829 && pixel_index <= 1830) || (pixel_index >= 1842 && pixel_index <= 1843) || (pixel_index >= 1854 && pixel_index <= 1856) || (pixel_index >= 1868 && pixel_index <= 1870) || (pixel_index >= 1880 && pixel_index <= 1881) || (pixel_index >= 1892 && pixel_index <= 1893) || (pixel_index >= 1905 && pixel_index <= 1907) || (pixel_index >= 1925 && pixel_index <= 1926) || (pixel_index >= 1938 && pixel_index <= 1939) || (pixel_index >= 1950 && pixel_index <= 1952) || (pixel_index >= 1964 && pixel_index <= 1966) || (pixel_index >= 1976 && pixel_index <= 1977) || (pixel_index >= 1988 && pixel_index <= 1989) || (pixel_index >= 2001 && pixel_index <= 2003) || (pixel_index >= 2021 && pixel_index <= 2022) || (pixel_index >= 2034 && pixel_index <= 2035) || (pixel_index >= 2046 && pixel_index <= 2048) || (pixel_index >= 2060 && pixel_index <= 2062) || (pixel_index >= 2072 && pixel_index <= 2073) || (pixel_index >= 2084 && pixel_index <= 2085) || (pixel_index >= 2097 && pixel_index <= 2099) || (pixel_index >= 2117 && pixel_index <= 2118) || (pixel_index >= 2130 && pixel_index <= 2132) || (pixel_index >= 2142 && pixel_index <= 2144) || (pixel_index >= 2156 && pixel_index <= 2158) || (pixel_index >= 2168 && pixel_index <= 2169) || (pixel_index >= 2180 && pixel_index <= 2181) || (pixel_index >= 2193 && pixel_index <= 2195) || (pixel_index >= 2213 && pixel_index <= 2214) || (pixel_index >= 2226 && pixel_index <= 2228) || (pixel_index >= 2238 && pixel_index <= 2240) || (pixel_index >= 2252 && pixel_index <= 2254) || (pixel_index >= 2264 && pixel_index <= 2265) || (pixel_index >= 2276 && pixel_index <= 2277) || (pixel_index >= 2289 && pixel_index <= 2291) || (pixel_index >= 2309 && pixel_index <= 2310) || (pixel_index >= 2334 && pixel_index <= 2336) || (pixel_index >= 2348 && pixel_index <= 2350) || (pixel_index >= 2360 && pixel_index <= 2361) || (pixel_index >= 2372 && pixel_index <= 2373) || (pixel_index >= 2385 && pixel_index <= 2387) || (pixel_index >= 2405 && pixel_index <= 2406) || (pixel_index >= 2430 && pixel_index <= 2432) || (pixel_index >= 2456 && pixel_index <= 2457) || (pixel_index >= 2468 && pixel_index <= 2469) || (pixel_index >= 2481 && pixel_index <= 2483) || (pixel_index >= 2501 && pixel_index <= 2502) || (pixel_index >= 2526 && pixel_index <= 2528) || (pixel_index >= 2552 && pixel_index <= 2553) || (pixel_index >= 2564 && pixel_index <= 2565) || (pixel_index >= 2577 && pixel_index <= 2579) || (pixel_index >= 2597 && pixel_index <= 2598) || (pixel_index >= 2606 && pixel_index <= 2607) || (pixel_index >= 2622 && pixel_index <= 2624) || (pixel_index >= 2648 && pixel_index <= 2649) || (pixel_index >= 2660 && pixel_index <= 2661) || (pixel_index >= 2673 && pixel_index <= 2675) || (pixel_index >= 2693 && pixel_index <= 2694) || (pixel_index >= 2702 && pixel_index <= 2703) || (pixel_index >= 2718 && pixel_index <= 2720) || (pixel_index >= 2744 && pixel_index <= 2745) || (pixel_index >= 2756 && pixel_index <= 2757) || (pixel_index >= 2769 && pixel_index <= 2771) || (pixel_index >= 2789 && pixel_index <= 2790) || (pixel_index >= 2798 && pixel_index <= 2799) || (pixel_index >= 2814 && pixel_index <= 2816) || (pixel_index >= 2840 && pixel_index <= 2841) || (pixel_index >= 2852 && pixel_index <= 2853) || (pixel_index >= 2865 && pixel_index <= 2867) || (pixel_index >= 2885 && pixel_index <= 2886) || (pixel_index >= 2894 && pixel_index <= 2895) || (pixel_index >= 2910 && pixel_index <= 2912) || (pixel_index >= 2924 && pixel_index <= 2926) || (pixel_index >= 2936 && pixel_index <= 2937) || (pixel_index >= 2948 && pixel_index <= 2949) || (pixel_index >= 2961 && pixel_index <= 2963) || (pixel_index >= 2981 && pixel_index <= 2982) || (pixel_index >= 2990 && pixel_index <= 2991) || (pixel_index >= 3006 && pixel_index <= 3008) || (pixel_index >= 3020 && pixel_index <= 3022) || (pixel_index >= 3032 && pixel_index <= 3033) || (pixel_index >= 3044 && pixel_index <= 3045) || (pixel_index >= 3057 && pixel_index <= 3059) || (pixel_index >= 3077 && pixel_index <= 3078) || (pixel_index >= 3090 && pixel_index <= 3091) || (pixel_index >= 3102 && pixel_index <= 3104) || (pixel_index >= 3116 && pixel_index <= 3118) || (pixel_index >= 3128 && pixel_index <= 3129) || (pixel_index >= 3140 && pixel_index <= 3141) || (pixel_index >= 3153 && pixel_index <= 3155) || (pixel_index >= 3173 && pixel_index <= 3174) || (pixel_index >= 3186 && pixel_index <= 3187) || (pixel_index >= 3198 && pixel_index <= 3200) || (pixel_index >= 3212 && pixel_index <= 3214) || (pixel_index >= 3224 && pixel_index <= 3225) || (pixel_index >= 3236 && pixel_index <= 3237) || (pixel_index >= 3249 && pixel_index <= 3251) || (pixel_index >= 3269 && pixel_index <= 3270) || (pixel_index >= 3282 && pixel_index <= 3283) || (pixel_index >= 3294 && pixel_index <= 3296) || (pixel_index >= 3308 && pixel_index <= 3310) || (pixel_index >= 3320 && pixel_index <= 3321) || (pixel_index >= 3332 && pixel_index <= 3333) || (pixel_index >= 3345 && pixel_index <= 3347) || (pixel_index >= 3365 && pixel_index <= 3366) || (pixel_index >= 3378 && pixel_index <= 3379) || (pixel_index >= 3390 && pixel_index <= 3392) || (pixel_index >= 3404 && pixel_index <= 3406) || (pixel_index >= 3416 && pixel_index <= 3417) || (pixel_index >= 3428 && pixel_index <= 3429) || (pixel_index >= 3441 && pixel_index <= 3443) || (pixel_index >= 3465 && pixel_index <= 3466) || (pixel_index >= 3486 && pixel_index <= 3488) || (pixel_index >= 3500 && pixel_index <= 3502) || (pixel_index >= 3512 && pixel_index <= 3513) || (pixel_index >= 3524 && pixel_index <= 3525) || (pixel_index >= 3561 && pixel_index <= 3562) || (pixel_index >= 3582 && pixel_index <= 3584) || (pixel_index >= 3596 && pixel_index <= 3598) || (pixel_index >= 3608 && pixel_index <= 3609) || (pixel_index >= 3620 && pixel_index <= 3621) || (pixel_index >= 3657 && pixel_index <= 3658) || (pixel_index >= 3678 && pixel_index <= 3680) || (pixel_index >= 3692 && pixel_index <= 3694) || (pixel_index >= 3704 && pixel_index <= 3705) || (pixel_index >= 3716 && pixel_index <= 3717) || (pixel_index >= 3753 && pixel_index <= 3754) || (pixel_index >= 3774 && pixel_index <= 3776) || (pixel_index >= 3788 && pixel_index <= 3790) || (pixel_index >= 3800 && pixel_index <= 3801) || (pixel_index >= 3812 && pixel_index <= 3813) || (pixel_index >= 3849 && pixel_index <= 3851) || (pixel_index >= 3870 && pixel_index <= 3872) || (pixel_index >= 3884 && pixel_index <= 3886) || (pixel_index >= 3896 && pixel_index <= 3898) || (pixel_index >= 3908 && pixel_index <= 3910)) begin
            oled_data = BLUE_HEX;
        end else if ((pixel_index >= 1356 && pixel_index <= 1364) || (pixel_index >= 1377 && pixel_index <= 1389) || (pixel_index >= 1403 && pixel_index <= 1406) || (pixel_index >= 1415 && pixel_index <= 1427) || (pixel_index >= 1451 && pixel_index <= 1460) || (pixel_index >= 1473 && pixel_index <= 1485) || (pixel_index >= 1498 && pixel_index <= 1502) || (pixel_index >= 1510 && pixel_index <= 1523) || (pixel_index >= 1547 && pixel_index <= 1556) || (pixel_index >= 1569 && pixel_index <= 1581) || (pixel_index >= 1594 && pixel_index <= 1598) || (pixel_index >= 1606 && pixel_index <= 1619) || (pixel_index >= 1643 && pixel_index <= 1652) || (pixel_index >= 1665 && pixel_index <= 1677) || (pixel_index >= 1690 && pixel_index <= 1694) || (pixel_index >= 1702 && pixel_index <= 1715) || (pixel_index >= 1740 && pixel_index <= 1748) || (pixel_index >= 1761 && pixel_index <= 1773) || (pixel_index >= 1786 && pixel_index <= 1790) || (pixel_index >= 1798 && pixel_index <= 1811) || (pixel_index >= 1831 && pixel_index <= 1835) || (pixel_index >= 1844 && pixel_index <= 1848) || (pixel_index >= 1857 && pixel_index <= 1860) || (pixel_index >= 1871 && pixel_index <= 1874) || (pixel_index >= 1882 && pixel_index <= 1886) || (pixel_index >= 1894 && pixel_index <= 1898) || (pixel_index >= 1908 && pixel_index <= 1912) || (pixel_index >= 1927 && pixel_index <= 1931) || (pixel_index >= 1940 && pixel_index <= 1944) || (pixel_index >= 1953 && pixel_index <= 1956) || (pixel_index >= 1967 && pixel_index <= 1970) || (pixel_index >= 1978 && pixel_index <= 1982) || (pixel_index >= 1990 && pixel_index <= 1994) || (pixel_index >= 2004 && pixel_index <= 2008) || (pixel_index >= 2023 && pixel_index <= 2027) || (pixel_index >= 2036 && pixel_index <= 2040) || (pixel_index >= 2049 && pixel_index <= 2052) || (pixel_index >= 2063 && pixel_index <= 2066) || (pixel_index >= 2074 && pixel_index <= 2078) || (pixel_index >= 2086 && pixel_index <= 2090) || (pixel_index >= 2100 && pixel_index <= 2104) || (pixel_index >= 2119 && pixel_index <= 2123) || (pixel_index >= 2133 && pixel_index <= 2136) || (pixel_index >= 2145 && pixel_index <= 2148) || (pixel_index >= 2159 && pixel_index <= 2162) || (pixel_index >= 2170 && pixel_index <= 2174) || (pixel_index >= 2182 && pixel_index <= 2186) || (pixel_index >= 2196 && pixel_index <= 2200) || (pixel_index >= 2215 && pixel_index <= 2219) || (pixel_index >= 2229 && pixel_index <= 2232) || (pixel_index >= 2241 && pixel_index <= 2244) || (pixel_index >= 2255 && pixel_index <= 2258) || (pixel_index >= 2266 && pixel_index <= 2270) || (pixel_index >= 2278 && pixel_index <= 2282) || (pixel_index >= 2292 && pixel_index <= 2296) || (pixel_index >= 2311 && pixel_index <= 2315) || (pixel_index >= 2337 && pixel_index <= 2340) || (pixel_index >= 2351 && pixel_index <= 2354) || (pixel_index >= 2362 && pixel_index <= 2366) || (pixel_index >= 2374 && pixel_index <= 2378) || (pixel_index >= 2388 && pixel_index <= 2392) || (pixel_index >= 2407 && pixel_index <= 2411) || (pixel_index >= 2433 && pixel_index <= 2450) || (pixel_index >= 2458 && pixel_index <= 2462) || (pixel_index >= 2470 && pixel_index <= 2474) || (pixel_index >= 2484 && pixel_index <= 2488) || (pixel_index >= 2503 && pixel_index <= 2507) || (pixel_index >= 2529 && pixel_index <= 2542) || (pixel_index >= 2554 && pixel_index <= 2558) || (pixel_index >= 2566 && pixel_index <= 2570) || (pixel_index >= 2580 && pixel_index <= 2584) || (pixel_index >= 2599 && pixel_index <= 2603) || (pixel_index >= 2608 && pixel_index <= 2616) || (pixel_index >= 2625 && pixel_index <= 2638) || (pixel_index >= 2650 && pixel_index <= 2654) || (pixel_index >= 2662 && pixel_index <= 2666) || (pixel_index >= 2676 && pixel_index <= 2680) || (pixel_index >= 2695 && pixel_index <= 2699) || (pixel_index >= 2704 && pixel_index <= 2712) || (pixel_index >= 2721 && pixel_index <= 2734) || (pixel_index >= 2746 && pixel_index <= 2750) || (pixel_index >= 2758 && pixel_index <= 2762) || (pixel_index >= 2772 && pixel_index <= 2776) || (pixel_index >= 2791 && pixel_index <= 2795) || (pixel_index >= 2800 && pixel_index <= 2808) || (pixel_index >= 2817 && pixel_index <= 2834) || (pixel_index >= 2842 && pixel_index <= 2846) || (pixel_index >= 2854 && pixel_index <= 2858) || (pixel_index >= 2868 && pixel_index <= 2872) || (pixel_index >= 2887 && pixel_index <= 2891) || (pixel_index >= 2896 && pixel_index <= 2904) || (pixel_index >= 2913 && pixel_index <= 2916) || (pixel_index >= 2927 && pixel_index <= 2930) || (pixel_index >= 2938 && pixel_index <= 2942) || (pixel_index >= 2950 && pixel_index <= 2954) || (pixel_index >= 2964 && pixel_index <= 2968) || (pixel_index >= 2983 && pixel_index <= 2987) || (pixel_index >= 2992 && pixel_index <= 3000) || (pixel_index >= 3009 && pixel_index <= 3012) || (pixel_index >= 3023 && pixel_index <= 3026) || (pixel_index >= 3034 && pixel_index <= 3038) || (pixel_index >= 3046 && pixel_index <= 3050) || (pixel_index >= 3060 && pixel_index <= 3064) || (pixel_index >= 3079 && pixel_index <= 3083) || (pixel_index >= 3092 && pixel_index <= 3096) || (pixel_index >= 3105 && pixel_index <= 3108) || (pixel_index >= 3119 && pixel_index <= 3122) || (pixel_index >= 3130 && pixel_index <= 3134) || (pixel_index >= 3142 && pixel_index <= 3146) || (pixel_index >= 3156 && pixel_index <= 3160) || (pixel_index >= 3175 && pixel_index <= 3179) || (pixel_index >= 3188 && pixel_index <= 3192) || (pixel_index >= 3201 && pixel_index <= 3204) || (pixel_index >= 3215 && pixel_index <= 3218) || (pixel_index >= 3226 && pixel_index <= 3230) || (pixel_index >= 3238 && pixel_index <= 3242) || (pixel_index >= 3252 && pixel_index <= 3256) || (pixel_index >= 3271 && pixel_index <= 3275) || (pixel_index >= 3284 && pixel_index <= 3288) || (pixel_index >= 3297 && pixel_index <= 3300) || (pixel_index >= 3311 && pixel_index <= 3314) || (pixel_index >= 3322 && pixel_index <= 3326) || (pixel_index >= 3334 && pixel_index <= 3338) || (pixel_index >= 3348 && pixel_index <= 3352) || (pixel_index >= 3367 && pixel_index <= 3371) || (pixel_index >= 3380 && pixel_index <= 3384) || (pixel_index >= 3393 && pixel_index <= 3396) || (pixel_index >= 3407 && pixel_index <= 3410) || (pixel_index >= 3418 && pixel_index <= 3422) || (pixel_index >= 3430 && pixel_index <= 3434) || (pixel_index >= 3444 && pixel_index <= 3448) || (pixel_index >= 3467 && pixel_index <= 3476) || (pixel_index >= 3489 && pixel_index <= 3492) || (pixel_index >= 3503 && pixel_index <= 3506) || (pixel_index >= 3514 && pixel_index <= 3518) || (pixel_index >= 3526 && pixel_index <= 3539) || (pixel_index >= 3563 && pixel_index <= 3572) || (pixel_index >= 3585 && pixel_index <= 3588) || (pixel_index >= 3599 && pixel_index <= 3602) || (pixel_index >= 3610 && pixel_index <= 3614) || (pixel_index >= 3622 && pixel_index <= 3635) || (pixel_index >= 3659 && pixel_index <= 3668) || (pixel_index >= 3681 && pixel_index <= 3684) || (pixel_index >= 3695 && pixel_index <= 3698) || (pixel_index >= 3706 && pixel_index <= 3710) || (pixel_index >= 3718 && pixel_index <= 3731) || (pixel_index >= 3755 && pixel_index <= 3764) || (pixel_index >= 3777 && pixel_index <= 3780) || (pixel_index >= 3791 && pixel_index <= 3794) || (pixel_index >= 3802 && pixel_index <= 3806) || (pixel_index >= 3814 && pixel_index <= 3827) || (pixel_index >= 3852 && pixel_index <= 3860) || (pixel_index >= 3873 && pixel_index <= 3876) || (pixel_index >= 3887 && pixel_index <= 3890) || (pixel_index >= 3899 && pixel_index <= 3902) || (pixel_index >= 3911 && pixel_index <= 3923) || (pixel_index >= 4136 && pixel_index <= 4138) || (pixel_index >= 4144 && pixel_index <= 4146) || (pixel_index >= 4152 && pixel_index <= 4155) || (pixel_index >= 4163 && pixel_index <= 4166) || (pixel_index >= 4173 && pixel_index <= 4180) || (pixel_index >= 4184 && pixel_index <= 4191) || (pixel_index >= 4195 && pixel_index <= 4201) || (pixel_index >= 4209 && pixel_index <= 4212) || (pixel_index >= 4232 && pixel_index <= 4234) || (pixel_index >= 4240 && pixel_index <= 4242) || (pixel_index >= 4248 && pixel_index <= 4251) || (pixel_index >= 4258 && pixel_index <= 4263) || (pixel_index >= 4269 && pixel_index <= 4276) || (pixel_index >= 4280 && pixel_index <= 4287) || (pixel_index >= 4291 && pixel_index <= 4297) || (pixel_index >= 4304 && pixel_index <= 4309) || (pixel_index >= 4328 && pixel_index <= 4332) || (pixel_index >= 4334 && pixel_index <= 4338) || (pixel_index >= 4342 && pixel_index <= 4343) || (pixel_index >= 4348 && pixel_index <= 4349) || (pixel_index >= 4353 && pixel_index <= 4354) || (pixel_index >= 4359 && pixel_index <= 4360) || (pixel_index >= 4368 && pixel_index <= 4369) || (pixel_index >= 4376 && pixel_index <= 4378) || (pixel_index >= 4387 && pixel_index <= 4389) || (pixel_index >= 4394 && pixel_index <= 4395) || (pixel_index >= 4399 && pixel_index <= 4400) || (pixel_index >= 4405 && pixel_index <= 4406) || (pixel_index >= 4424 && pixel_index <= 4428) || (pixel_index >= 4430 && pixel_index <= 4434) || (pixel_index >= 4438 && pixel_index <= 4439) || (pixel_index >= 4444 && pixel_index <= 4445) || (pixel_index >= 4449 && pixel_index <= 4450) || (pixel_index >= 4455 && pixel_index <= 4456) || (pixel_index >= 4464 && pixel_index <= 4465) || (pixel_index >= 4472 && pixel_index <= 4474) || (pixel_index >= 4483 && pixel_index <= 4485) || (pixel_index >= 4490 && pixel_index <= 4491) || (pixel_index >= 4495 && pixel_index <= 4496) || (pixel_index >= 4501 && pixel_index <= 4502) || (pixel_index >= 4520 && pixel_index <= 4522) || (pixel_index >= 4524 && pixel_index <= 4526) || (pixel_index >= 4528 && pixel_index <= 4530) || (pixel_index >= 4534 && pixel_index <= 4535) || (pixel_index >= 4540 && pixel_index <= 4541) || (pixel_index >= 4545 && pixel_index <= 4546) || (pixel_index >= 4560 && pixel_index <= 4561) || (pixel_index >= 4568 && pixel_index <= 4570) || (pixel_index >= 4579 && pixel_index <= 4581) || (pixel_index >= 4586 && pixel_index <= 4587) || (pixel_index >= 4591 && pixel_index <= 4592) || (pixel_index >= 4616 && pixel_index <= 4618) || (pixel_index >= 4620 && pixel_index <= 4622) || (pixel_index >= 4624 && pixel_index <= 4626) || (pixel_index >= 4630 && pixel_index <= 4637) || (pixel_index >= 4643 && pixel_index <= 4646) || (pixel_index >= 4656 && pixel_index <= 4657) || (pixel_index >= 4664 && pixel_index <= 4669) || (pixel_index >= 4675 && pixel_index <= 4682) || (pixel_index >= 4689 && pixel_index <= 4692) || (pixel_index >= 4712 && pixel_index <= 4714) || (pixel_index >= 4720 && pixel_index <= 4722) || (pixel_index >= 4726 && pixel_index <= 4733) || (pixel_index >= 4740 && pixel_index <= 4744) || (pixel_index >= 4752 && pixel_index <= 4753) || (pixel_index >= 4760 && pixel_index <= 4765) || (pixel_index >= 4771 && pixel_index <= 4778) || (pixel_index >= 4786 && pixel_index <= 4790) || (pixel_index >= 4808 && pixel_index <= 4810) || (pixel_index >= 4816 && pixel_index <= 4818) || (pixel_index >= 4822 && pixel_index <= 4823) || (pixel_index >= 4828 && pixel_index <= 4829) || (pixel_index >= 4833 && pixel_index <= 4834) || (pixel_index >= 4839 && pixel_index <= 4840) || (pixel_index >= 4848 && pixel_index <= 4849) || (pixel_index >= 4856 && pixel_index <= 4858) || (pixel_index >= 4867 && pixel_index <= 4869) || (pixel_index >= 4874 && pixel_index <= 4875) || (pixel_index >= 4879 && pixel_index <= 4880) || (pixel_index >= 4885 && pixel_index <= 4886) || (pixel_index >= 4904 && pixel_index <= 4906) || (pixel_index >= 4912 && pixel_index <= 4914) || (pixel_index >= 4918 && pixel_index <= 4919) || (pixel_index >= 4924 && pixel_index <= 4925) || (pixel_index >= 4929 && pixel_index <= 4930) || (pixel_index >= 4935 && pixel_index <= 4936) || (pixel_index >= 4944 && pixel_index <= 4945) || (pixel_index >= 4952 && pixel_index <= 4954) || (pixel_index >= 4963 && pixel_index <= 4965) || (pixel_index >= 4970 && pixel_index <= 4971) || (pixel_index >= 4975 && pixel_index <= 4976) || (pixel_index >= 4981 && pixel_index <= 4982) || (pixel_index >= 5000 && pixel_index <= 5002) || (pixel_index >= 5008 && pixel_index <= 5010) || (pixel_index >= 5014 && pixel_index <= 5015) || (pixel_index >= 5020 && pixel_index <= 5021) || (pixel_index >= 5025 && pixel_index <= 5032) || (pixel_index >= 5040 && pixel_index <= 5041) || (pixel_index >= 5048 && pixel_index <= 5055) || (pixel_index >= 5059 && pixel_index <= 5061) || (pixel_index >= 5066 && pixel_index <= 5067) || (pixel_index >= 5071 && pixel_index <= 5078) || (pixel_index >= 5096 && pixel_index <= 5098) || (pixel_index >= 5104 && pixel_index <= 5106) || (pixel_index >= 5110 && pixel_index <= 5111) || (pixel_index >= 5116 && pixel_index <= 5117) || (pixel_index >= 5123 && pixel_index <= 5126) || (pixel_index >= 5136 && pixel_index <= 5137) || (pixel_index >= 5144 && pixel_index <= 5151) || (pixel_index >= 5155 && pixel_index <= 5157) || (pixel_index >= 5162 && pixel_index <= 5163) || (pixel_index >= 5169 && pixel_index <= 5172)) begin
            oled_data = WHITE_HEX;
        end else begin
            oled_data = BG_BLUE_HEX;
        end
    end
endmodule
